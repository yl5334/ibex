

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO mult8x8 
  PIN a[7] 
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.7719 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 101.123 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END a[7]
  PIN a[6] 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.622 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.9649 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.237 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END a[6]
  PIN a[5] 
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.1404 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 91.386 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END a[5]
  PIN a[4] 
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.2807 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.105 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END a[4]
  PIN a[3] 
    ANTENNAPARTIALMETALAREA 2.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.362 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.6491 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 104.368 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END a[3]
  PIN a[2] 
    ANTENNAPARTIALMETALAREA 1.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.5789 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.0088 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END a[2]
  PIN a[1] 
    ANTENNAPARTIALMETALAREA 2.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.474 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.6491 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 104.368 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END a[1]
  PIN a[0] 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.622 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.2105 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 102.746 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END a[0]
  PIN b[7] 
    ANTENNAPARTIALMETALAREA 2.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.4035 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.86 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END b[7]
  PIN b[6] 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.3333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 99.5 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END b[6]
  PIN b[5] 
    ANTENNAPARTIALMETALAREA 2.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.362 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.1579 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 117.351 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END b[5]
  PIN b[4] 
    ANTENNAPARTIALMETALAREA 1.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.4561 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 96.2544 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END b[4]
  PIN b[3] 
    ANTENNAPARTIALMETALAREA 2.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.474 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.3468 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 107.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END b[3]
  PIN b[2] 
    ANTENNAPARTIALMETALAREA 1.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.7018 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 89.7632 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END b[2]
  PIN b[1] 
    ANTENNAPARTIALMETALAREA 1.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.586 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.2632 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 88.1404 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END b[1]
  PIN b[0] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.806 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.9825 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 135.202 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL ;
  END b[0]
  PIN result[15] 
    ANTENNAPARTIALMETALAREA 2.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.026 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.66 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.01389 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.80198 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.024024 LAYER VL ;
  END result[15]
  PIN result[14] 
    ANTENNAPARTIALMETALAREA 4.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.242 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.603 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.07576 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.7841 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0461007 LAYER VL ;
  END result[14]
  PIN result[13] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.602 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.49716 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.63213 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0461184 LAYER VL ;
  END result[13]
  PIN result[12] 
    ANTENNAPARTIALMETALAREA 3.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.47 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.603 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.58402 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.9078 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0461007 LAYER VL ;
  END result[12]
  PIN result[11] 
    ANTENNAPARTIALMETALAREA 3.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.986 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.602 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.71238 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 6.42844 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0461184 LAYER VL ;
  END result[11]
  PIN result[10] 
    ANTENNAPARTIALMETALAREA 3.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.174 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.603 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.46108 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.45294 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0461007 LAYER VL ;
  END result[10]
  PIN result[9] 
    ANTENNAPARTIALMETALAREA 3.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.766 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.603 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.46108 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.45294 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0461007 LAYER VL ;
  END result[9]
  PIN result[8] 
    ANTENNAPARTIALMETALAREA 2.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.99 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.602 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.29731 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.8927 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0461184 LAYER VL ;
  END result[8]
  PIN result[7] 
    ANTENNAPARTIALMETALAREA 4.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.058 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.602 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.11207 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.9073 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0461184 LAYER VL ;
  END result[7]
  PIN result[6] 
    ANTENNAPARTIALMETALAREA 3.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.358 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.893 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.21046 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.03212 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0845219 LAYER VL ;
  END result[6]
  PIN result[5] 
    ANTENNAPARTIALMETALAREA 4.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.058 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.893 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.78098 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 10.1431 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0845219 LAYER VL ;
  END result[5]
  PIN result[4] 
    ANTENNAPARTIALMETALAREA 4.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.466 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.848 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.94747 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.14466 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0561798 LAYER VL ;
  END result[4]
  PIN result[3] 
    ANTENNAPARTIALMETALAREA 6.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.346 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.014 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.91976 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 14.6616 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0794439 LAYER VL ;
  END result[3]
  PIN result[2] 
    ANTENNAPARTIALMETALAREA 5.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.386 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.014 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.6854 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.9168 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0794439 LAYER VL ;
  END result[2]
  PIN result[1] 
    ANTENNAPARTIALMETALAREA 5.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.314 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.014 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.67349 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 14.03 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0794439 LAYER VL ;
  END result[1]
  PIN result[0] 
    ANTENNAPARTIALMETALAREA 6.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.458 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.014 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.78073 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 14.1472 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0794439 LAYER VL ;
  END result[0]
  PIN clk 
    ANTENNAPARTIALMETALAREA 10.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 37.666 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5544 LAYER M2 ; 
    ANTENNAMAXAREACAR 20.5931 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 77.728 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER V2 ;
    ANTENNAMAXCUTCAR 1.22655 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 132.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 498.464 LAYER M3 ;
    ANTENNAGATEAREA 28.9728 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.1712 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 94.9325 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.52525 LAYER VL ;
  END clk
  PIN resetn 
    ANTENNAPARTIALMETALAREA 1.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.204 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.9451 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 36.9275 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.196078 LAYER V2 ;
  END resetn
END mult8x8

END LIBRARY
