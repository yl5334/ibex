

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO ibex_top 
  PIN clk_i 
    ANTENNAPARTIALMETALAREA 1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 62.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 234.432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5976 LAYER M3 ; 
    ANTENNAMAXAREACAR 151.904 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 575.449 LAYER M3 ;
    ANTENNAMAXCUTCAR 5.55556 LAYER VL ;
  END clk_i
  PIN rst_ni 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.7703 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END rst_ni
  PIN test_en_i 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.3739 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 116.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END test_en_i
  PIN ram_cfg_i[9] 
  END ram_cfg_i[9]
  PIN ram_cfg_i[8] 
  END ram_cfg_i[8]
  PIN ram_cfg_i[7] 
  END ram_cfg_i[7]
  PIN ram_cfg_i[6] 
  END ram_cfg_i[6]
  PIN ram_cfg_i[5] 
  END ram_cfg_i[5]
  PIN ram_cfg_i[4] 
  END ram_cfg_i[4]
  PIN ram_cfg_i[3] 
  END ram_cfg_i[3]
  PIN ram_cfg_i[2] 
  END ram_cfg_i[2]
  PIN ram_cfg_i[1] 
  END ram_cfg_i[1]
  PIN ram_cfg_i[0] 
  END ram_cfg_i[0]
  PIN hart_id_i[31] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.9685 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 96.3559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[31]
  PIN hart_id_i[30] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 42.1892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[30]
  PIN hart_id_i[29] 
    ANTENNAPARTIALMETALAREA 4.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.096 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 48.3919 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 183.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[29]
  PIN hart_id_i[28] 
    ANTENNAPARTIALMETALAREA 2.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.62 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.7252 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 121.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[28]
  PIN hart_id_i[27] 
    ANTENNAPARTIALMETALAREA 2.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.1757 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 123.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[27]
  PIN hart_id_i[26] 
    ANTENNAPARTIALMETALAREA 3.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.284 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.8333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 151.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[26]
  PIN hart_id_i[25] 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.3739 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 116.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[25]
  PIN hart_id_i[24] 
    ANTENNAPARTIALMETALAREA 2.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.436 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.0225 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 111.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[24]
  PIN hart_id_i[23] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.5721 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[23]
  PIN hart_id_i[22] 
    ANTENNAPARTIALMETALAREA 2.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.732 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.527 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 128.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[22]
  PIN hart_id_i[21] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.8694 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 99.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[21]
  PIN hart_id_i[20] 
    ANTENNAPARTIALMETALAREA 2.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.324 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.8243 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 118.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[20]
  PIN hart_id_i[19] 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.7703 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[19]
  PIN hart_id_i[18] 
    ANTENNAPARTIALMETALAREA 3.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.654 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.9144 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 175.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[18]
  PIN hart_id_i[17] 
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.7703 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[17]
  PIN hart_id_i[16] 
    ANTENNAPARTIALMETALAREA 2.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.732 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.9234 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[16]
  PIN hart_id_i[15] 
    ANTENNAPARTIALMETALAREA 2.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.5721 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[15]
  PIN hart_id_i[14] 
    ANTENNAPARTIALMETALAREA 2.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.212 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.2297 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 138.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[14]
  PIN hart_id_i[13] 
    ANTENNAPARTIALMETALAREA 2.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.473 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 113.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[13]
  PIN hart_id_i[12] 
    ANTENNAPARTIALMETALAREA 3.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.506 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 43.6622 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 163.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[12]
  PIN hart_id_i[11] 
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.9775 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 129.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[11]
  PIN hart_id_i[10] 
    ANTENNAPARTIALMETALAREA 2.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.62 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.6261 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 124.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[10]
  PIN hart_id_i[9] 
    ANTENNAPARTIALMETALAREA 2.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.7793 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 136.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[9]
  PIN hart_id_i[8] 
    ANTENNAPARTIALMETALAREA 4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.948 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 48.8423 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 184.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[8]
  PIN hart_id_i[7] 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.8694 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 99.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[7]
  PIN hart_id_i[6] 
    ANTENNAPARTIALMETALAREA 2.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.804 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.536 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 161.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[6]
  PIN hart_id_i[5] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.806 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.5991 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 115.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[5]
  PIN hart_id_i[4] 
    ANTENNAPARTIALMETALAREA 2.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.212 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.2297 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 138.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[4]
  PIN hart_id_i[3] 
    ANTENNAPARTIALMETALAREA 1.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.0766 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 126.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[3]
  PIN hart_id_i[2] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.07658 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 35.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[2]
  PIN hart_id_i[1] 
    ANTENNAPARTIALMETALAREA 2.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.2748 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 119.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[1]
  PIN hart_id_i[0] 
    ANTENNAPARTIALMETALAREA 2.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.732 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.6892 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 174.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[0]
  PIN boot_addr_i[31] 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.812 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.65315 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 38.0225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[31]
  PIN boot_addr_i[30] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.4459 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 105.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[30]
  PIN boot_addr_i[29] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[29]
  PIN boot_addr_i[28] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.6441 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 98.8559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[28]
  PIN boot_addr_i[27] 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.812 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.65315 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 38.0225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[27]
  PIN boot_addr_i[26] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[26]
  PIN boot_addr_i[25] 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.812 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.65315 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 38.0225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[25]
  PIN boot_addr_i[24] 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.516 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.95045 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 29.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[24]
  PIN boot_addr_i[23] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.6441 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 98.8559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[23]
  PIN boot_addr_i[22] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.3468 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 108.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[22]
  PIN boot_addr_i[21] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.6712 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 106.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[21]
  PIN boot_addr_i[20] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.4459 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 105.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[20]
  PIN boot_addr_i[19] 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.516 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 8.75225 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 34.6892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[19]
  PIN boot_addr_i[18] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.545 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 102.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[18]
  PIN boot_addr_i[17] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[17]
  PIN boot_addr_i[16] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.3739 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 116.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[16]
  PIN boot_addr_i[15] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.0766 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 126.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[15]
  PIN boot_addr_i[14] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.7793 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 136.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[14]
  PIN boot_addr_i[13] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.2748 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 119.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[13]
  PIN boot_addr_i[12] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.1757 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 123.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[12]
  PIN boot_addr_i[11] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.0766 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 126.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[11]
  PIN boot_addr_i[10] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.36 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.8784 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 133.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[10]
  PIN boot_addr_i[9] 
    ANTENNAPARTIALMETALAREA 0.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 8.97748 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 37.1892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[9]
  PIN boot_addr_i[8] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.7793 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 136.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[8]
  PIN boot_addr_i[7] 
  END boot_addr_i[7]
  PIN boot_addr_i[6] 
  END boot_addr_i[6]
  PIN boot_addr_i[5] 
  END boot_addr_i[5]
  PIN boot_addr_i[4] 
  END boot_addr_i[4]
  PIN boot_addr_i[3] 
  END boot_addr_i[3]
  PIN boot_addr_i[2] 
  END boot_addr_i[2]
  PIN boot_addr_i[1] 
  END boot_addr_i[1]
  PIN boot_addr_i[0] 
  END boot_addr_i[0]
  PIN instr_req_o 
    ANTENNAPARTIALMETALAREA 3.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.284 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4672 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.8799 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 21.6086 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.11111 LAYER VL ;
  END instr_req_o
  PIN instr_gnt_i 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.258 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.5991 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 117.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_gnt_i
  PIN instr_rvalid_i 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.0946 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 100.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rvalid_i
  PIN instr_addr_o[31] 
    ANTENNAPARTIALMETALAREA 8.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.708 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.88445 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 10.8057 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[31]
  PIN instr_addr_o[30] 
    ANTENNAPARTIALMETALAREA 6.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.42 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.10581 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.82562 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END instr_addr_o[30]
  PIN instr_addr_o[29] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.252 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.790282 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.00069 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[29]
  PIN instr_addr_o[28] 
    ANTENNAPARTIALMETALAREA 4.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.5 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.47 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.6089 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[28]
  PIN instr_addr_o[27] 
    ANTENNAPARTIALMETALAREA 1.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.476 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.806899 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.0184 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[27]
  PIN instr_addr_o[26] 
    ANTENNAPARTIALMETALAREA 1.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.66 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.35309 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.74599 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END instr_addr_o[26]
  PIN instr_addr_o[25] 
    ANTENNAPARTIALMETALAREA 1.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.476 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.696909 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2.61622 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[25]
  PIN instr_addr_o[24] 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.62 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.39998 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.32186 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END instr_addr_o[24]
  PIN instr_addr_o[23] 
    ANTENNAPARTIALMETALAREA 1.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.476 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.93865 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.50712 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END instr_addr_o[23]
  PIN instr_addr_o[22] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.86842 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 6.95321 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[22]
  PIN instr_addr_o[21] 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.812 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.461103 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.72957 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[21]
  PIN instr_addr_o[20] 
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.3794 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.10485 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[20]
  PIN instr_addr_o[19] 
    ANTENNAPARTIALMETALAREA 3.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.06 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.28089 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.89189 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END instr_addr_o[19]
  PIN instr_addr_o[18] 
    ANTENNAPARTIALMETALAREA 1.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.18 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.946958 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.55331 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END instr_addr_o[18]
  PIN instr_addr_o[17] 
    ANTENNAPARTIALMETALAREA 0.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.404 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.560015 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2.09555 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[17]
  PIN instr_addr_o[16] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.44923 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.04906 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[16]
  PIN instr_addr_o[15] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.252 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.935485 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.53076 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[15]
  PIN instr_addr_o[14] 
    ANTENNAPARTIALMETALAREA 1.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.548 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.928759 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.50712 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END instr_addr_o[14]
  PIN instr_addr_o[13] 
    ANTENNAPARTIALMETALAREA 1.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.996 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.661696 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2.48239 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END instr_addr_o[13]
  PIN instr_addr_o[12] 
    ANTENNAPARTIALMETALAREA 4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.244 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.4253 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.39832 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END instr_addr_o[12]
  PIN instr_addr_o[11] 
    ANTENNAPARTIALMETALAREA 3.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.876 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.20294 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.58417 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[11]
  PIN instr_addr_o[10] 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.844 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.88959 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.35153 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END instr_addr_o[10]
  PIN instr_addr_o[9] 
    ANTENNAPARTIALMETALAREA 2.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.916 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.07436 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.07181 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[9]
  PIN instr_addr_o[8] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.90344 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 10.7383 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END instr_addr_o[8]
  PIN instr_addr_o[7] 
    ANTENNAPARTIALMETALAREA 5.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.572 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.84468 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.01454 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END instr_addr_o[7]
  PIN instr_addr_o[6] 
    ANTENNAPARTIALMETALAREA 5.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.98 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.64805 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 6.26766 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[6]
  PIN instr_addr_o[5] 
    ANTENNAPARTIALMETALAREA 0.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.965158 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.60396 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[5]
  PIN instr_addr_o[4] 
    ANTENNAPARTIALMETALAREA 1.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.772 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.899085 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.36073 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END instr_addr_o[4]
  PIN instr_addr_o[3] 
    ANTENNAPARTIALMETALAREA 0.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.768521 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2.90376 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END instr_addr_o[3]
  PIN instr_addr_o[2] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.886424 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.26667 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0296736 LAYER VL ;
  END instr_addr_o[2]
  PIN instr_rdata_i[31] 
    ANTENNAPARTIALMETALAREA 1.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.218 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.536 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 70.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[31]
  PIN instr_rdata_i[30] 
    ANTENNAPARTIALMETALAREA 0.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.554 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.8964 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 107.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[30]
  PIN instr_rdata_i[29] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.258 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.3468 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[29]
  PIN instr_rdata_i[28] 
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.146 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.5 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 120.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[28]
  PIN instr_rdata_i[27] 
    ANTENNAPARTIALMETALAREA 0.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.626 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.8333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 60.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[27]
  PIN instr_rdata_i[26] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.258 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.9955 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[26]
  PIN instr_rdata_i[25] 
    ANTENNAPARTIALMETALAREA 0.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.2027 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 130.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[25]
  PIN instr_rdata_i[24] 
    ANTENNAPARTIALMETALAREA 0.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.554 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.7973 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[24]
  PIN instr_rdata_i[23] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.33 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.1306 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 50.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[23]
  PIN instr_rdata_i[22] 
    ANTENNAPARTIALMETALAREA 0.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.922 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.9324 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 57.1892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[22]
  PIN instr_rdata_i[21] 
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.146 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.5991 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 117.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[21]
  PIN instr_rdata_i[20] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.8964 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 107.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[20]
  PIN instr_rdata_i[19] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.258 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.9955 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[19]
  PIN instr_rdata_i[18] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.258 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.9955 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[18]
  PIN instr_rdata_i[17] 
    ANTENNAPARTIALMETALAREA 2.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.844 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.3198 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 101.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[17]
  PIN instr_rdata_i[16] 
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.146 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.6982 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 113.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[16]
  PIN instr_rdata_i[15] 
    ANTENNAPARTIALMETALAREA 0.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.1036 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 133.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[15]
  PIN instr_rdata_i[14] 
    ANTENNAPARTIALMETALAREA 1.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.514 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.4369 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 73.8559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[14]
  PIN instr_rdata_i[13] 
    ANTENNAPARTIALMETALAREA 0.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.5 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 120.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[13]
  PIN instr_rdata_i[12] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.258 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.9955 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[12]
  PIN instr_rdata_i[11] 
    ANTENNAPARTIALMETALAREA 2.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.3468 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[11]
  PIN instr_rdata_i[10] 
    ANTENNAPARTIALMETALAREA 0.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.7523 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 130.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[10]
  PIN instr_rdata_i[9] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.8694 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 98.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[9]
  PIN instr_rdata_i[8] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.6982 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 113.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[8]
  PIN instr_rdata_i[7] 
    ANTENNAPARTIALMETALAREA 0.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.554 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.8964 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 107.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[7]
  PIN instr_rdata_i[6] 
    ANTENNAPARTIALMETALAREA 0.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.3018 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 127.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[6]
  PIN instr_rdata_i[5] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.5811 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 141.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[5]
  PIN instr_rdata_i[4] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.7072 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 147.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[4]
  PIN instr_rdata_i[3] 
    ANTENNAPARTIALMETALAREA 0.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.5 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 120.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[3]
  PIN instr_rdata_i[2] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.8964 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 107.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[2]
  PIN instr_rdata_i[1] 
    ANTENNAPARTIALMETALAREA 2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.548 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.0225 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 111.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[1]
  PIN instr_rdata_i[0] 
    ANTENNAPARTIALMETALAREA 1.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.8423 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.8559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[0]
  PIN instr_rdata_intg_i[6] 
  END instr_rdata_intg_i[6]
  PIN instr_rdata_intg_i[5] 
  END instr_rdata_intg_i[5]
  PIN instr_rdata_intg_i[4] 
  END instr_rdata_intg_i[4]
  PIN instr_rdata_intg_i[3] 
  END instr_rdata_intg_i[3]
  PIN instr_rdata_intg_i[2] 
  END instr_rdata_intg_i[2]
  PIN instr_rdata_intg_i[1] 
  END instr_rdata_intg_i[1]
  PIN instr_rdata_intg_i[0] 
  END instr_rdata_intg_i[0]
  PIN instr_err_i 
    ANTENNAPARTIALMETALAREA 1.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.218 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.1396 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 83.8559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_err_i
  PIN data_req_o 
    ANTENNAPARTIALMETALAREA 0.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.182 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.64 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.3314 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 42.25 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.25 LAYER VL ;
  END data_req_o
  PIN data_gnt_i 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 29.0225 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 109.689 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_gnt_i
  PIN data_rvalid_i 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 24.518 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 93.0225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rvalid_i
  PIN data_we_o 
    ANTENNAPARTIALMETALAREA 6.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.754 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.9224 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.1019 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 150.801 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.68817 LAYER VL ;
  END data_we_o
  PIN data_be_o[3] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.592 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.63596 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 6.09753 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0617284 LAYER VL ;
  END data_be_o[3]
  PIN data_be_o[2] 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.698 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.92 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.968323 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.61691 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0395648 LAYER VL ;
  END data_be_o[2]
  PIN data_be_o[1] 
    ANTENNAPARTIALMETALAREA 2.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.286 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.01877 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.73907 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0197824 LAYER V2 ;
  END data_be_o[1]
  PIN data_be_o[0] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.16 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.78 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 10.2838 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.137931 LAYER VL ;
  END data_be_o[0]
  PIN data_addr_o[31] 
    ANTENNAPARTIALMETALAREA 30.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 114.404 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 33.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 126.984 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.0236 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.2364 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 79.8677 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END data_addr_o[31]
  PIN data_addr_o[30] 
    ANTENNAPARTIALMETALAREA 5.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.61 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 79.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 298.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.0236 LAYER M3 ; 
    ANTENNAMAXAREACAR 63.1109 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 240.584 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_addr_o[30]
  PIN data_addr_o[29] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 107.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 401.08 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0828 LAYER M3 ; 
    ANTENNAMAXAREACAR 72.1554 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 271.376 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.77305 LAYER VL ;
  END data_addr_o[29]
  PIN data_addr_o[28] 
    ANTENNAPARTIALMETALAREA 4.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.058 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 107.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 407.296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1964 LAYER M3 ; 
    ANTENNAMAXAREACAR 60.1203 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 232.306 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END data_addr_o[28]
  PIN data_addr_o[27] 
    ANTENNAPARTIALMETALAREA 22.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 84.286 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 29.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 113.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.0956 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.7622 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 60.0734 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.746269 LAYER VL ;
  END data_addr_o[27]
  PIN data_addr_o[26] 
    ANTENNAPARTIALMETALAREA 38.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 143.042 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 139.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 518.296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.0236 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.9208 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 149.289 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_addr_o[26]
  PIN data_addr_o[25] 
    ANTENNAPARTIALMETALAREA 27.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 101.898 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 124.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 462.352 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.0956 LAYER M3 ; 
    ANTENNAMAXAREACAR 72.1251 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 268.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END data_addr_o[25]
  PIN data_addr_o[24] 
    ANTENNAPARTIALMETALAREA 14.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 54.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 55.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 207.496 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.0236 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.4565 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 107.748 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_addr_o[24]
  PIN data_addr_o[23] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 78.736 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6328 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.0685 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 120.961 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.41844 LAYER VL ;
  END data_addr_o[23]
  PIN data_addr_o[22] 
    ANTENNAPARTIALMETALAREA 4.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.982 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 75.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 283.272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 60.7009 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 242.006 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END data_addr_o[22]
  PIN data_addr_o[21] 
    ANTENNAPARTIALMETALAREA 57.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 213.046 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 51.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 192.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2556 LAYER M3 ; 
    ANTENNAMAXAREACAR 97.8747 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 373.654 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.77305 LAYER VL ;
  END data_addr_o[21]
  PIN data_addr_o[20] 
    ANTENNAPARTIALMETALAREA 63.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 234.358 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 42.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 157.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.4448 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 85.9151 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END data_addr_o[20]
  PIN data_addr_o[19] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 45.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 170.496 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.6355 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 112.002 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END data_addr_o[19]
  PIN data_addr_o[18] 
    ANTENNAPARTIALMETALAREA 63.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 234.654 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 76.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 289.192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1964 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.1026 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 188.384 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END data_addr_o[18]
  PIN data_addr_o[17] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 59.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 220.52 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.21 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.9591 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 127.325 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.78571 LAYER VL ;
  END data_addr_o[17]
  PIN data_addr_o[16] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 99.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 373.552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1964 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.56 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 138.706 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END data_addr_o[16]
  PIN data_addr_o[15] 
    ANTENNAPARTIALMETALAREA 1.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.734 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 86.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 323.232 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.4472 LAYER M3 ; 
    ANTENNAMAXAREACAR 88.5676 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 334.754 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END data_addr_o[15]
  PIN data_addr_o[14] 
    ANTENNAPARTIALMETALAREA 29.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 108.854 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 81.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 306.656 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2556 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.2607 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 197.548 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END data_addr_o[14]
  PIN data_addr_o[13] 
    ANTENNAPARTIALMETALAREA 1.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 44.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 170.792 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2844 LAYER M3 ; 
    ANTENNAMAXAREACAR 120.695 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 451.415 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.38095 LAYER VL ;
  END data_addr_o[13]
  PIN data_addr_o[12] 
    ANTENNAPARTIALMETALAREA 2.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.99 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 41.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 155.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.21 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.4294 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 138.111 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.97619 LAYER VL ;
  END data_addr_o[12]
  PIN data_addr_o[11] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.47 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 44.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 172.272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.978 LAYER M3 ; 
    ANTENNAMAXAREACAR 62.8624 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 243.032 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.97619 LAYER VL ;
  END data_addr_o[11]
  PIN data_addr_o[10] 
    ANTENNAPARTIALMETALAREA 3.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.95 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 70.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 266.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.905 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.9025 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END data_addr_o[10]
  PIN data_addr_o[9] 
    ANTENNAPARTIALMETALAREA 5.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.83 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 97.384 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0372 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.2424 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 55.5995 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.78571 LAYER VL ;
  END data_addr_o[9]
  PIN data_addr_o[8] 
    ANTENNAPARTIALMETALAREA 16.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 62.086 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 76.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 290.376 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.4472 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.7246 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 139.418 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.68817 LAYER VL ;
  END data_addr_o[8]
  PIN data_addr_o[7] 
    ANTENNAPARTIALMETALAREA 18.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 69.19 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 74.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 278.536 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.4472 LAYER M3 ; 
    ANTENNAMAXAREACAR 48.0411 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 183.671 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.68817 LAYER VL ;
  END data_addr_o[7]
  PIN data_addr_o[6] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.51 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 97.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 368.52 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.4472 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.241 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 510.314 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END data_addr_o[6]
  PIN data_addr_o[5] 
    ANTENNAPARTIALMETALAREA 4.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.686 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 76.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 286.232 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4572 LAYER M3 ; 
    ANTENNAMAXAREACAR 68.2321 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 259.876 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.38095 LAYER VL ;
  END data_addr_o[5]
  PIN data_addr_o[4] 
    ANTENNAPARTIALMETALAREA 47.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 174.714 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4572 LAYER M3 ; 
    ANTENNAMAXAREACAR 73.8706 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 284.467 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.68817 LAYER VL ;
  END data_addr_o[4]
  PIN data_addr_o[3] 
    ANTENNAPARTIALMETALAREA 16.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.346 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 61.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 233.544 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2844 LAYER M3 ; 
    ANTENNAMAXAREACAR 49.4801 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 190.583 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.38095 LAYER VL ;
  END data_addr_o[3]
  PIN data_addr_o[2] 
    ANTENNAPARTIALMETALAREA 5.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.942 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 50.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 188.848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3156 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.0534 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.474 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END data_addr_o[2]
  PIN data_wdata_o[31] 
    ANTENNAPARTIALMETALAREA 3.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.67386 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 6.19792 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0189394 LAYER V2 ;
  END data_wdata_o[31]
  PIN data_wdata_o[30] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.18409 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.40417 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[30]
  PIN data_wdata_o[29] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.47 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.6928 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 6.26799 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0189394 LAYER V2 ;
  END data_wdata_o[29]
  PIN data_wdata_o[28] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.55076 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.88258 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[28]
  PIN data_wdata_o[27] 
    ANTENNAPARTIALMETALAREA 3.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.766 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.056 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.16061 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 11.7689 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[27]
  PIN data_wdata_o[26] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.51 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.41439 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 20.178 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[26]
  PIN data_wdata_o[25] 
    ANTENNAPARTIALMETALAREA 3.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.174 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.568 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.4447 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.0303 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[25]
  PIN data_wdata_o[24] 
    ANTENNAPARTIALMETALAREA 5.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.534 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.92 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.27424 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.83182 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[24]
  PIN data_wdata_o[23] 
    ANTENNAPARTIALMETALAREA 4.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.022 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.25038 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 8.34261 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER V2 ;
  END data_wdata_o[23]
  PIN data_wdata_o[22] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.344 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.65758 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 32.3095 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[22]
  PIN data_wdata_o[21] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.68 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.48712 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 35.5254 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[21]
  PIN data_wdata_o[20] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.69848 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.9417 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[20]
  PIN data_wdata_o[19] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.208 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.11894 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.98485 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[19]
  PIN data_wdata_o[18] 
    ANTENNAPARTIALMETALAREA 4.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.318 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.96629 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 15.6949 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER V2 ;
  END data_wdata_o[18]
  PIN data_wdata_o[17] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.15682 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.125 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[17]
  PIN data_wdata_o[16] 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.214 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 77.256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.4076 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 38.9913 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[16]
  PIN data_wdata_o[15] 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.142 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 72.52 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.7402 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 43.5833 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[15]
  PIN data_wdata_o[14] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.99091 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 11.3095 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[14]
  PIN data_wdata_o[13] 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 102.712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.8318 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 55.2375 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[13]
  PIN data_wdata_o[12] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.214 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 78.736 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.3386 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 38.3977 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[12]
  PIN data_wdata_o[11] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.784 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.80833 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 17.9356 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[11]
  PIN data_wdata_o[10] 
    ANTENNAPARTIALMETALAREA 3.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.766 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.344 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.08182 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 15.3057 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[10]
  PIN data_wdata_o[9] 
    ANTENNAPARTIALMETALAREA 6.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.086 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.963636 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.64015 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[9]
  PIN data_wdata_o[8] 
    ANTENNAPARTIALMETALAREA 3.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.95 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 94.424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.4606 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 46.3473 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[8]
  PIN data_wdata_o[7] 
    ANTENNAPARTIALMETALAREA 3.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.874 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.512 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.09621 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.20076 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[7]
  PIN data_wdata_o[6] 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.698 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 38.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 143.56 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.6341 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 69.0909 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[6]
  PIN data_wdata_o[5] 
    ANTENNAPARTIALMETALAREA 4.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.466 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.20417 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 8.16004 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0189394 LAYER V2 ;
  END data_wdata_o[5]
  PIN data_wdata_o[4] 
    ANTENNAPARTIALMETALAREA 4.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.686 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 101.232 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.4076 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 49.711 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[4]
  PIN data_wdata_o[3] 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.698 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 74 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.0205 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 37.453 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[3]
  PIN data_wdata_o[2] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 29.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 110.704 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.7402 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 62.0833 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[2]
  PIN data_wdata_o[1] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.576 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.89545 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 29.5682 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[1]
  PIN data_wdata_o[0] 
    ANTENNAPARTIALMETALAREA 6.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.53182 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 24.2424 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[0]
  PIN data_rdata_i[31] 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.844 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 24.518 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 94.6892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[31]
  PIN data_rdata_i[30] 
    ANTENNAPARTIALMETALAREA 3.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.504 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 45.2387 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 169.689 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[30]
  PIN data_rdata_i[29] 
    ANTENNAPARTIALMETALAREA 1.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.846 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.0586 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 59.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[29]
  PIN data_rdata_i[28] 
    ANTENNAPARTIALMETALAREA 1.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.75225 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 36.3559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[28]
  PIN data_rdata_i[27] 
    ANTENNAPARTIALMETALAREA 2.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 26.3198 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 99.6892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[27]
  PIN data_rdata_i[26] 
    ANTENNAPARTIALMETALAREA 1.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.846 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.6712 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 106.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[26]
  PIN data_rdata_i[25] 
    ANTENNAPARTIALMETALAREA 2.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.102 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 28.7973 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 108.856 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[25]
  PIN data_rdata_i[24] 
    ANTENNAPARTIALMETALAREA 2.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 27.2207 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[24]
  PIN data_rdata_i[23] 
    ANTENNAPARTIALMETALAREA 1.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 23.6171 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 89.6892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[23]
  PIN data_rdata_i[22] 
    ANTENNAPARTIALMETALAREA 2.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 25.4189 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 96.3559 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[22]
  PIN data_rdata_i[21] 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 29.0225 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 109.689 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[21]
  PIN data_rdata_i[20] 
    ANTENNAPARTIALMETALAREA 0.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.182 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.6171 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[20]
  PIN data_rdata_i[19] 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.698 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.6171 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[19]
  PIN data_rdata_i[18] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.328 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.2748 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 119.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[18]
  PIN data_rdata_i[17] 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 24.518 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 93.0225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[17]
  PIN data_rdata_i[16] 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.622 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.8604 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 66.3559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[16]
  PIN data_rdata_i[15] 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 24.518 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 93.0225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[15]
  PIN data_rdata_i[14] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.1667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 89.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[14]
  PIN data_rdata_i[13] 
    ANTENNAPARTIALMETALAREA 1.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.6622 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 73.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[13]
  PIN data_rdata_i[12] 
    ANTENNAPARTIALMETALAREA 0.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.182 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.9685 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 96.3559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[12]
  PIN data_rdata_i[11] 
    ANTENNAPARTIALMETALAREA 0.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.182 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.464 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 79.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[11]
  PIN data_rdata_i[10] 
    ANTENNAPARTIALMETALAREA 1.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.85135 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 33.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[10]
  PIN data_rdata_i[9] 
    ANTENNAPARTIALMETALAREA 2.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 27.2207 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[9]
  PIN data_rdata_i[8] 
    ANTENNAPARTIALMETALAREA 2.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 25.4189 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 96.3559 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[8]
  PIN data_rdata_i[7] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.5721 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[7]
  PIN data_rdata_i[6] 
    ANTENNAPARTIALMETALAREA 2.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 28.1216 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 106.356 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[6]
  PIN data_rdata_i[5] 
    ANTENNAPARTIALMETALAREA 1.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 23.6171 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 89.6892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[5]
  PIN data_rdata_i[4] 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.698 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.3739 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 116.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[4]
  PIN data_rdata_i[3] 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 24.518 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 93.0225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[3]
  PIN data_rdata_i[2] 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.142 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.5541 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 43.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[2]
  PIN data_rdata_i[1] 
    ANTENNAPARTIALMETALAREA 2.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.99 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.3559 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 49.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[1]
  PIN data_rdata_i[0] 
    ANTENNAPARTIALMETALAREA 0.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.182 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.7703 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[0]
  PIN data_rdata_intg_i[6] 
  END data_rdata_intg_i[6]
  PIN data_rdata_intg_i[5] 
  END data_rdata_intg_i[5]
  PIN data_rdata_intg_i[4] 
  END data_rdata_intg_i[4]
  PIN data_rdata_intg_i[3] 
  END data_rdata_intg_i[3]
  PIN data_rdata_intg_i[2] 
  END data_rdata_intg_i[2]
  PIN data_rdata_intg_i[1] 
  END data_rdata_intg_i[1]
  PIN data_rdata_intg_i[0] 
  END data_rdata_intg_i[0]
  PIN data_err_i 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 24.518 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 93.0225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_err_i
  PIN irq_software_i 
    ANTENNAPARTIALMETALAREA 2.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.62 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.6261 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 124.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_software_i
  PIN irq_timer_i 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.7703 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_timer_i
  PIN irq_external_i 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.7793 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 45.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_external_i
  PIN irq_fast_i[14] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.5721 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[14]
  PIN irq_fast_i[13] 
    ANTENNAPARTIALMETALAREA 2.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.99 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.1577 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 148.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[13]
  PIN irq_fast_i[12] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.8694 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 99.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[12]
  PIN irq_fast_i[11] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.694 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.8063 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 145.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[11]
  PIN irq_fast_i[10] 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.994 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.1396 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 83.8559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[10]
  PIN irq_fast_i[9] 
    ANTENNAPARTIALMETALAREA 2.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.842 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.8063 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 143.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[9]
  PIN irq_fast_i[8] 
    ANTENNAPARTIALMETALAREA 2.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.7523 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 130.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[8]
  PIN irq_fast_i[7] 
    ANTENNAPARTIALMETALAREA 2.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.732 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.8333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 151.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[7]
  PIN irq_fast_i[6] 
    ANTENNAPARTIALMETALAREA 1.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.7703 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[6]
  PIN irq_fast_i[5] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.694 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.3018 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 128.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[5]
  PIN irq_fast_i[4] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.3378 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 77.1892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[4]
  PIN irq_fast_i[3] 
    ANTENNAPARTIALMETALAREA 0.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.59 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.7793 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 45.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[3]
  PIN irq_fast_i[2] 
    ANTENNAPARTIALMETALAREA 2.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.1757 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 123.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[2]
  PIN irq_fast_i[1] 
    ANTENNAPARTIALMETALAREA 0.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.59 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.7793 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 45.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[1]
  PIN irq_fast_i[0] 
    ANTENNAPARTIALMETALAREA 2.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.1 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.6802 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 141.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[0]
  PIN irq_nm_i 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.214 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.7973 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 108.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_nm_i
  PIN scramble_key_valid_i 
  END scramble_key_valid_i
  PIN scramble_key_i[127] 
  END scramble_key_i[127]
  PIN scramble_key_i[126] 
  END scramble_key_i[126]
  PIN scramble_key_i[125] 
  END scramble_key_i[125]
  PIN scramble_key_i[124] 
  END scramble_key_i[124]
  PIN scramble_key_i[123] 
  END scramble_key_i[123]
  PIN scramble_key_i[122] 
  END scramble_key_i[122]
  PIN scramble_key_i[121] 
  END scramble_key_i[121]
  PIN scramble_key_i[120] 
  END scramble_key_i[120]
  PIN scramble_key_i[119] 
  END scramble_key_i[119]
  PIN scramble_key_i[118] 
  END scramble_key_i[118]
  PIN scramble_key_i[117] 
  END scramble_key_i[117]
  PIN scramble_key_i[116] 
  END scramble_key_i[116]
  PIN scramble_key_i[115] 
  END scramble_key_i[115]
  PIN scramble_key_i[114] 
  END scramble_key_i[114]
  PIN scramble_key_i[113] 
  END scramble_key_i[113]
  PIN scramble_key_i[112] 
  END scramble_key_i[112]
  PIN scramble_key_i[111] 
  END scramble_key_i[111]
  PIN scramble_key_i[110] 
  END scramble_key_i[110]
  PIN scramble_key_i[109] 
  END scramble_key_i[109]
  PIN scramble_key_i[108] 
  END scramble_key_i[108]
  PIN scramble_key_i[107] 
  END scramble_key_i[107]
  PIN scramble_key_i[106] 
  END scramble_key_i[106]
  PIN scramble_key_i[105] 
  END scramble_key_i[105]
  PIN scramble_key_i[104] 
  END scramble_key_i[104]
  PIN scramble_key_i[103] 
  END scramble_key_i[103]
  PIN scramble_key_i[102] 
  END scramble_key_i[102]
  PIN scramble_key_i[101] 
  END scramble_key_i[101]
  PIN scramble_key_i[100] 
  END scramble_key_i[100]
  PIN scramble_key_i[99] 
  END scramble_key_i[99]
  PIN scramble_key_i[98] 
  END scramble_key_i[98]
  PIN scramble_key_i[97] 
  END scramble_key_i[97]
  PIN scramble_key_i[96] 
  END scramble_key_i[96]
  PIN scramble_key_i[95] 
  END scramble_key_i[95]
  PIN scramble_key_i[94] 
  END scramble_key_i[94]
  PIN scramble_key_i[93] 
  END scramble_key_i[93]
  PIN scramble_key_i[92] 
  END scramble_key_i[92]
  PIN scramble_key_i[91] 
  END scramble_key_i[91]
  PIN scramble_key_i[90] 
  END scramble_key_i[90]
  PIN scramble_key_i[89] 
  END scramble_key_i[89]
  PIN scramble_key_i[88] 
  END scramble_key_i[88]
  PIN scramble_key_i[87] 
  END scramble_key_i[87]
  PIN scramble_key_i[86] 
  END scramble_key_i[86]
  PIN scramble_key_i[85] 
  END scramble_key_i[85]
  PIN scramble_key_i[84] 
  END scramble_key_i[84]
  PIN scramble_key_i[83] 
  END scramble_key_i[83]
  PIN scramble_key_i[82] 
  END scramble_key_i[82]
  PIN scramble_key_i[81] 
  END scramble_key_i[81]
  PIN scramble_key_i[80] 
  END scramble_key_i[80]
  PIN scramble_key_i[79] 
  END scramble_key_i[79]
  PIN scramble_key_i[78] 
  END scramble_key_i[78]
  PIN scramble_key_i[77] 
  END scramble_key_i[77]
  PIN scramble_key_i[76] 
  END scramble_key_i[76]
  PIN scramble_key_i[75] 
  END scramble_key_i[75]
  PIN scramble_key_i[74] 
  END scramble_key_i[74]
  PIN scramble_key_i[73] 
  END scramble_key_i[73]
  PIN scramble_key_i[72] 
  END scramble_key_i[72]
  PIN scramble_key_i[71] 
  END scramble_key_i[71]
  PIN scramble_key_i[70] 
  END scramble_key_i[70]
  PIN scramble_key_i[69] 
  END scramble_key_i[69]
  PIN scramble_key_i[68] 
  END scramble_key_i[68]
  PIN scramble_key_i[67] 
  END scramble_key_i[67]
  PIN scramble_key_i[66] 
  END scramble_key_i[66]
  PIN scramble_key_i[65] 
  END scramble_key_i[65]
  PIN scramble_key_i[64] 
  END scramble_key_i[64]
  PIN scramble_key_i[63] 
  END scramble_key_i[63]
  PIN scramble_key_i[62] 
  END scramble_key_i[62]
  PIN scramble_key_i[61] 
  END scramble_key_i[61]
  PIN scramble_key_i[60] 
  END scramble_key_i[60]
  PIN scramble_key_i[59] 
  END scramble_key_i[59]
  PIN scramble_key_i[58] 
  END scramble_key_i[58]
  PIN scramble_key_i[57] 
  END scramble_key_i[57]
  PIN scramble_key_i[56] 
  END scramble_key_i[56]
  PIN scramble_key_i[55] 
  END scramble_key_i[55]
  PIN scramble_key_i[54] 
  END scramble_key_i[54]
  PIN scramble_key_i[53] 
  END scramble_key_i[53]
  PIN scramble_key_i[52] 
  END scramble_key_i[52]
  PIN scramble_key_i[51] 
  END scramble_key_i[51]
  PIN scramble_key_i[50] 
  END scramble_key_i[50]
  PIN scramble_key_i[49] 
  END scramble_key_i[49]
  PIN scramble_key_i[48] 
  END scramble_key_i[48]
  PIN scramble_key_i[47] 
  END scramble_key_i[47]
  PIN scramble_key_i[46] 
  END scramble_key_i[46]
  PIN scramble_key_i[45] 
  END scramble_key_i[45]
  PIN scramble_key_i[44] 
  END scramble_key_i[44]
  PIN scramble_key_i[43] 
  END scramble_key_i[43]
  PIN scramble_key_i[42] 
  END scramble_key_i[42]
  PIN scramble_key_i[41] 
  END scramble_key_i[41]
  PIN scramble_key_i[40] 
  END scramble_key_i[40]
  PIN scramble_key_i[39] 
  END scramble_key_i[39]
  PIN scramble_key_i[38] 
  END scramble_key_i[38]
  PIN scramble_key_i[37] 
  END scramble_key_i[37]
  PIN scramble_key_i[36] 
  END scramble_key_i[36]
  PIN scramble_key_i[35] 
  END scramble_key_i[35]
  PIN scramble_key_i[34] 
  END scramble_key_i[34]
  PIN scramble_key_i[33] 
  END scramble_key_i[33]
  PIN scramble_key_i[32] 
  END scramble_key_i[32]
  PIN scramble_key_i[31] 
  END scramble_key_i[31]
  PIN scramble_key_i[30] 
  END scramble_key_i[30]
  PIN scramble_key_i[29] 
  END scramble_key_i[29]
  PIN scramble_key_i[28] 
  END scramble_key_i[28]
  PIN scramble_key_i[27] 
  END scramble_key_i[27]
  PIN scramble_key_i[26] 
  END scramble_key_i[26]
  PIN scramble_key_i[25] 
  END scramble_key_i[25]
  PIN scramble_key_i[24] 
  END scramble_key_i[24]
  PIN scramble_key_i[23] 
  END scramble_key_i[23]
  PIN scramble_key_i[22] 
  END scramble_key_i[22]
  PIN scramble_key_i[21] 
  END scramble_key_i[21]
  PIN scramble_key_i[20] 
  END scramble_key_i[20]
  PIN scramble_key_i[19] 
  END scramble_key_i[19]
  PIN scramble_key_i[18] 
  END scramble_key_i[18]
  PIN scramble_key_i[17] 
  END scramble_key_i[17]
  PIN scramble_key_i[16] 
  END scramble_key_i[16]
  PIN scramble_key_i[15] 
  END scramble_key_i[15]
  PIN scramble_key_i[14] 
  END scramble_key_i[14]
  PIN scramble_key_i[13] 
  END scramble_key_i[13]
  PIN scramble_key_i[12] 
  END scramble_key_i[12]
  PIN scramble_key_i[11] 
  END scramble_key_i[11]
  PIN scramble_key_i[10] 
  END scramble_key_i[10]
  PIN scramble_key_i[9] 
  END scramble_key_i[9]
  PIN scramble_key_i[8] 
  END scramble_key_i[8]
  PIN scramble_key_i[7] 
  END scramble_key_i[7]
  PIN scramble_key_i[6] 
  END scramble_key_i[6]
  PIN scramble_key_i[5] 
  END scramble_key_i[5]
  PIN scramble_key_i[4] 
  END scramble_key_i[4]
  PIN scramble_key_i[3] 
  END scramble_key_i[3]
  PIN scramble_key_i[2] 
  END scramble_key_i[2]
  PIN scramble_key_i[1] 
  END scramble_key_i[1]
  PIN scramble_key_i[0] 
  END scramble_key_i[0]
  PIN scramble_nonce_i[63] 
  END scramble_nonce_i[63]
  PIN scramble_nonce_i[62] 
  END scramble_nonce_i[62]
  PIN scramble_nonce_i[61] 
  END scramble_nonce_i[61]
  PIN scramble_nonce_i[60] 
  END scramble_nonce_i[60]
  PIN scramble_nonce_i[59] 
  END scramble_nonce_i[59]
  PIN scramble_nonce_i[58] 
  END scramble_nonce_i[58]
  PIN scramble_nonce_i[57] 
  END scramble_nonce_i[57]
  PIN scramble_nonce_i[56] 
  END scramble_nonce_i[56]
  PIN scramble_nonce_i[55] 
  END scramble_nonce_i[55]
  PIN scramble_nonce_i[54] 
  END scramble_nonce_i[54]
  PIN scramble_nonce_i[53] 
  END scramble_nonce_i[53]
  PIN scramble_nonce_i[52] 
  END scramble_nonce_i[52]
  PIN scramble_nonce_i[51] 
  END scramble_nonce_i[51]
  PIN scramble_nonce_i[50] 
  END scramble_nonce_i[50]
  PIN scramble_nonce_i[49] 
  END scramble_nonce_i[49]
  PIN scramble_nonce_i[48] 
  END scramble_nonce_i[48]
  PIN scramble_nonce_i[47] 
  END scramble_nonce_i[47]
  PIN scramble_nonce_i[46] 
  END scramble_nonce_i[46]
  PIN scramble_nonce_i[45] 
  END scramble_nonce_i[45]
  PIN scramble_nonce_i[44] 
  END scramble_nonce_i[44]
  PIN scramble_nonce_i[43] 
  END scramble_nonce_i[43]
  PIN scramble_nonce_i[42] 
  END scramble_nonce_i[42]
  PIN scramble_nonce_i[41] 
  END scramble_nonce_i[41]
  PIN scramble_nonce_i[40] 
  END scramble_nonce_i[40]
  PIN scramble_nonce_i[39] 
  END scramble_nonce_i[39]
  PIN scramble_nonce_i[38] 
  END scramble_nonce_i[38]
  PIN scramble_nonce_i[37] 
  END scramble_nonce_i[37]
  PIN scramble_nonce_i[36] 
  END scramble_nonce_i[36]
  PIN scramble_nonce_i[35] 
  END scramble_nonce_i[35]
  PIN scramble_nonce_i[34] 
  END scramble_nonce_i[34]
  PIN scramble_nonce_i[33] 
  END scramble_nonce_i[33]
  PIN scramble_nonce_i[32] 
  END scramble_nonce_i[32]
  PIN scramble_nonce_i[31] 
  END scramble_nonce_i[31]
  PIN scramble_nonce_i[30] 
  END scramble_nonce_i[30]
  PIN scramble_nonce_i[29] 
  END scramble_nonce_i[29]
  PIN scramble_nonce_i[28] 
  END scramble_nonce_i[28]
  PIN scramble_nonce_i[27] 
  END scramble_nonce_i[27]
  PIN scramble_nonce_i[26] 
  END scramble_nonce_i[26]
  PIN scramble_nonce_i[25] 
  END scramble_nonce_i[25]
  PIN scramble_nonce_i[24] 
  END scramble_nonce_i[24]
  PIN scramble_nonce_i[23] 
  END scramble_nonce_i[23]
  PIN scramble_nonce_i[22] 
  END scramble_nonce_i[22]
  PIN scramble_nonce_i[21] 
  END scramble_nonce_i[21]
  PIN scramble_nonce_i[20] 
  END scramble_nonce_i[20]
  PIN scramble_nonce_i[19] 
  END scramble_nonce_i[19]
  PIN scramble_nonce_i[18] 
  END scramble_nonce_i[18]
  PIN scramble_nonce_i[17] 
  END scramble_nonce_i[17]
  PIN scramble_nonce_i[16] 
  END scramble_nonce_i[16]
  PIN scramble_nonce_i[15] 
  END scramble_nonce_i[15]
  PIN scramble_nonce_i[14] 
  END scramble_nonce_i[14]
  PIN scramble_nonce_i[13] 
  END scramble_nonce_i[13]
  PIN scramble_nonce_i[12] 
  END scramble_nonce_i[12]
  PIN scramble_nonce_i[11] 
  END scramble_nonce_i[11]
  PIN scramble_nonce_i[10] 
  END scramble_nonce_i[10]
  PIN scramble_nonce_i[9] 
  END scramble_nonce_i[9]
  PIN scramble_nonce_i[8] 
  END scramble_nonce_i[8]
  PIN scramble_nonce_i[7] 
  END scramble_nonce_i[7]
  PIN scramble_nonce_i[6] 
  END scramble_nonce_i[6]
  PIN scramble_nonce_i[5] 
  END scramble_nonce_i[5]
  PIN scramble_nonce_i[4] 
  END scramble_nonce_i[4]
  PIN scramble_nonce_i[3] 
  END scramble_nonce_i[3]
  PIN scramble_nonce_i[2] 
  END scramble_nonce_i[2]
  PIN scramble_nonce_i[1] 
  END scramble_nonce_i[1]
  PIN scramble_nonce_i[0] 
  END scramble_nonce_i[0]
  PIN debug_req_i 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.7703 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END debug_req_i
  PIN crash_dump_o[159] 
    ANTENNAPARTIALMETALAREA 8.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.488 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 57.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 217.56 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5676 LAYER M3 ; 
    ANTENNAMAXAREACAR 57.2137 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 219.701 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.01149 LAYER VL ;
  END crash_dump_o[159]
  PIN crash_dump_o[158] 
    ANTENNAPARTIALMETALAREA 14.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 54.908 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.52 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4432 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.5423 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 154.872 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[158]
  PIN crash_dump_o[157] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 100.936 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.412 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.9989 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 117.57 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.84615 LAYER VL ;
  END crash_dump_o[157]
  PIN crash_dump_o[156] 
    ANTENNAPARTIALMETALAREA 13.84 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 51.652 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.848 LAYER M2 ; 
    ANTENNAMAXAREACAR 5.22605 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 19.4447 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0842697 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER M3 ;
    ANTENNAGATEAREA 3.4432 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.8721 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 76.0662 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.39578 LAYER VL ;
  END crash_dump_o[156]
  PIN crash_dump_o[155] 
    ANTENNAPARTIALMETALAREA 12.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 46.472 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.848 LAYER M2 ; 
    ANTENNAMAXAREACAR 5.21482 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 19.5742 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0842697 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 64.232 LAYER M3 ;
    ANTENNAGATEAREA 3.412 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.6601 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 49.8894 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.5641 LAYER VL ;
  END crash_dump_o[155]
  PIN crash_dump_o[154] 
    ANTENNAPARTIALMETALAREA 4.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.54 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4432 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.2173 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 97.7999 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[154]
  PIN crash_dump_o[153] 
    ANTENNAPARTIALMETALAREA 4.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.872 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.848 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.82718 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 6.75506 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0842697 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.88 LAYER M3 ;
    ANTENNAGATEAREA 3.412 LAYER M3 ; 
    ANTENNAMAXAREACAR 41.572 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 154.576 LAYER M3 ;
    ANTENNAMAXCUTCAR 5.12821 LAYER VL ;
  END crash_dump_o[153]
  PIN crash_dump_o[152] 
    ANTENNAPARTIALMETALAREA 8.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.044 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.848 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.03055 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 11.1556 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0561798 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.232 LAYER M3 ;
    ANTENNAGATEAREA 3.4432 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.1607 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 60.0756 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[152]
  PIN crash_dump_o[151] 
    ANTENNAPARTIALMETALAREA 0.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2972 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.8206 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 79.471 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[151]
  PIN crash_dump_o[150] 
    ANTENNAPARTIALMETALAREA 3.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.468 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.448 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2756 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.5919 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 67.7211 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER VL ;
  END crash_dump_o[150]
  PIN crash_dump_o[149] 
    ANTENNAPARTIALMETALAREA 0.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 31.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 120.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.412 LAYER M3 ; 
    ANTENNAMAXAREACAR 64.3222 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 242.409 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.62037 LAYER VL ;
  END crash_dump_o[149]
  PIN crash_dump_o[148] 
    ANTENNAPARTIALMETALAREA 1.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.996 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.014 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.98893 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 7.93664 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.119166 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 96.792 LAYER M3 ;
    ANTENNAGATEAREA 2.2156 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.4474 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 72.8497 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[148]
  PIN crash_dump_o[147] 
    ANTENNAPARTIALMETALAREA 5.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.904 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.014 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.86142 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 14.6203 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0794439 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.08 LAYER M3 ;
    ANTENNAGATEAREA 2.2756 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.5616 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 60.0138 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[147]
  PIN crash_dump_o[146] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2156 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.9676 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 85.8746 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[146]
  PIN crash_dump_o[145] 
    ANTENNAPARTIALMETALAREA 0.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 101.824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2156 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.8847 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 102.314 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER VL ;
  END crash_dump_o[145]
  PIN crash_dump_o[144] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.336 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4432 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.2266 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 65.5008 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.39578 LAYER VL ;
  END crash_dump_o[144]
  PIN crash_dump_o[143] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 44.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 167.536 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2968 LAYER M3 ; 
    ANTENNAMAXAREACAR 108.667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 417.908 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.84615 LAYER VL ;
  END crash_dump_o[143]
  PIN crash_dump_o[142] 
    ANTENNAPARTIALMETALAREA 1.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.66 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 42.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 160.432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3928 LAYER M3 ; 
    ANTENNAMAXAREACAR 62.5087 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 239.144 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.77305 LAYER VL ;
  END crash_dump_o[142]
  PIN crash_dump_o[141] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 53.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 202.464 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3568 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.9883 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 157.367 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.77225 LAYER VL ;
  END crash_dump_o[141]
  PIN crash_dump_o[140] 
    ANTENNAPARTIALMETALAREA 2.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.14 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 57.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 214.304 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5512 LAYER M3 ; 
    ANTENNAMAXAREACAR 52.8428 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 197.573 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[140]
  PIN crash_dump_o[139] 
    ANTENNAPARTIALMETALAREA 0.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 103.6 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2756 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.8269 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 65.2156 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[139]
  PIN crash_dump_o[138] 
    ANTENNAPARTIALMETALAREA 0.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 35.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 134.68 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1936 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.4123 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 88.3408 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[138]
  PIN crash_dump_o[137] 
    ANTENNAPARTIALMETALAREA 1.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.736 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.014 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.18039 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 8.69573 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.119166 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 98.272 LAYER M3 ;
    ANTENNAGATEAREA 2.2756 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.0791 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 87.6411 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[137]
  PIN crash_dump_o[136] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 46.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 174.344 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1312 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.2834 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 85.3688 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER VL ;
  END crash_dump_o[136]
  PIN crash_dump_o[135] 
    ANTENNAPARTIALMETALAREA 6.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.384 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 30.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 113.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2756 LAYER M3 ; 
    ANTENNAMAXAREACAR 55.3744 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 212.841 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[135]
  PIN crash_dump_o[134] 
    ANTENNAPARTIALMETALAREA 1.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.18 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 93.536 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.848 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.771 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 36.4685 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0561798 LAYER VL ;
  END crash_dump_o[134]
  PIN crash_dump_o[133] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 40.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 151.256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1096 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.6319 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 192.449 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[133]
  PIN crash_dump_o[132] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 134.088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1096 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.3078 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 116.448 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.768773 LAYER VL ;
  END crash_dump_o[132]
  PIN crash_dump_o[131] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 38.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 145.928 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1096 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.2342 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 131.528 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END crash_dump_o[131]
  PIN crash_dump_o[130] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 29.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 110.112 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.848 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.962 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 40.6652 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0561798 LAYER VL ;
  END crash_dump_o[130]
  PIN crash_dump_o[129] 
    ANTENNAPARTIALMETALAREA 0.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.96 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 71.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 266.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4044 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.6755 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 125.489 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[129]
  PIN crash_dump_o[127] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 30.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 111.888 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.5588 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.7327 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 82.5189 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[127]
  PIN crash_dump_o[126] 
    ANTENNAPARTIALMETALAREA 1.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.772 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 91.168 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0544 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.407 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 105.036 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[126]
  PIN crash_dump_o[125] 
    ANTENNAPARTIALMETALAREA 0.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 77.848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6812 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.8831 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.5 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[125]
  PIN crash_dump_o[124] 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.516 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1648 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.5348 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 150.135 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[124]
  PIN crash_dump_o[123] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6812 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.9974 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 49.2835 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.955763 LAYER VL ;
  END crash_dump_o[123]
  PIN crash_dump_o[122] 
    ANTENNAPARTIALMETALAREA 1.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.66 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0544 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.62322 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 32.2423 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[122]
  PIN crash_dump_o[121] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6812 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.6953 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 59.7191 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[121]
  PIN crash_dump_o[120] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1648 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.5738 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 59.7693 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.17391 LAYER VL ;
  END crash_dump_o[120]
  PIN crash_dump_o[119] 
    ANTENNAPARTIALMETALAREA 1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.784 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6812 LAYER M3 ; 
    ANTENNAMAXAREACAR 61.9594 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 235.697 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[119]
  PIN crash_dump_o[118] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.608 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1648 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.5235 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 57.734 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[118]
  PIN crash_dump_o[117] 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 89.984 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6812 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.0654 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 115.86 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[117]
  PIN crash_dump_o[116] 
    ANTENNAPARTIALMETALAREA 0.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.404 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 92.944 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1648 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.2404 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 57.2276 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[116]
  PIN crash_dump_o[115] 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 86.432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6812 LAYER M3 ; 
    ANTENNAMAXAREACAR 52.9706 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 199.924 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[115]
  PIN crash_dump_o[114] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 80.512 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1648 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.6302 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 102.414 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[114]
  PIN crash_dump_o[113] 
    ANTENNAPARTIALMETALAREA 0.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 88.208 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5152 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.1778 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 101.149 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[113]
  PIN crash_dump_o[112] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.896 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1648 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.0849 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 70.6306 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[112]
  PIN crash_dump_o[111] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 119.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6812 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.8655 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 156.16 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.86111 LAYER VL ;
  END crash_dump_o[111]
  PIN crash_dump_o[110] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 104.192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1648 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.9242 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 77.6028 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[110]
  PIN crash_dump_o[109] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 37.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 138.232 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6812 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.538 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 115.947 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[109]
  PIN crash_dump_o[108] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 29 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 108.04 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0544 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.998 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 59.1705 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[108]
  PIN crash_dump_o[107] 
    ANTENNAPARTIALMETALAREA 2.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.174 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 35.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 134.088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5152 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.7424 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 158.407 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.77778 LAYER VL ;
  END crash_dump_o[107]
  PIN crash_dump_o[106] 
    ANTENNAPARTIALMETALAREA 0.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 101.824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1648 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.5677 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 122 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.77778 LAYER VL ;
  END crash_dump_o[106]
  PIN crash_dump_o[105] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 102.416 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0784 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.5886 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 100.633 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[105]
  PIN crash_dump_o[104] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 121.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1648 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.5454 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 70.0782 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[104]
  PIN crash_dump_o[103] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 55.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 204.536 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6812 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.7514 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 126.954 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[103]
  PIN crash_dump_o[102] 
    ANTENNAPARTIALMETALAREA 1.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.996 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 120.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1648 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.5062 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 72.0491 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[102]
  PIN crash_dump_o[101] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 39.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 149.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1696 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.5729 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 117.116 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[101]
  PIN crash_dump_o[100] 
    ANTENNAPARTIALMETALAREA 1.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.292 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 34.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 127.28 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.554 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.6008 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 77.8321 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[100]
  PIN crash_dump_o[99] 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 36.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 137.048 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1048 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.581 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 84.6671 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[99]
  PIN crash_dump_o[98] 
    ANTENNAPARTIALMETALAREA 1.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.292 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 74.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 278.24 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4336 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.5866 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 135.666 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[98]
  PIN crash_dump_o[97] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 106.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 396.936 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3804 LAYER M3 ; 
    ANTENNAMAXAREACAR 77.2331 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 295.388 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[97]
  PIN crash_dump_o[95] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 131.128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.4474 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 50.6606 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[95]
  PIN crash_dump_o[94] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 30.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 113.96 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.5566 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 58.0395 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[94]
  PIN crash_dump_o[93] 
    ANTENNAPARTIALMETALAREA 1.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 94.72 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.20915 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 31.8383 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[93]
  PIN crash_dump_o[92] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 95.016 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.1796 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 38.1047 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[92]
  PIN crash_dump_o[91] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.896 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.19025 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 27.7258 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[91]
  PIN crash_dump_o[90] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.788 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.0564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 101.535 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[90]
  PIN crash_dump_o[89] 
    ANTENNAPARTIALMETALAREA 4.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.28 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 78.736 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.3761 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 48.0441 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER VL ;
  END crash_dump_o[89]
  PIN crash_dump_o[88] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 99.16 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.644 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 86.9783 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.77305 LAYER VL ;
  END crash_dump_o[88]
  PIN crash_dump_o[87] 
    ANTENNAPARTIALMETALAREA 1.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.504 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.7163 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 95.3908 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[87]
  PIN crash_dump_o[86] 
    ANTENNAPARTIALMETALAREA 2.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.916 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 28.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 105.968 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.8101 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 81.9336 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02881 LAYER VL ;
  END crash_dump_o[86]
  PIN crash_dump_o[85] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 36.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 138.824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.5505 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 120.333 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[85]
  PIN crash_dump_o[84] 
    ANTENNAPARTIALMETALAREA 0.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.404 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 34.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 130.832 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.0848 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.2228 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.77305 LAYER VL ;
  END crash_dump_o[84]
  PIN crash_dump_o[83] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 91.168 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.3026 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 59.1832 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.77305 LAYER VL ;
  END crash_dump_o[83]
  PIN crash_dump_o[82] 
    ANTENNAPARTIALMETALAREA 1.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.66 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 89.688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.0459 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 155.34 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.77305 LAYER VL ;
  END crash_dump_o[82]
  PIN crash_dump_o[81] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 33.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 128.464 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.2536 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 134.586 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.77305 LAYER VL ;
  END crash_dump_o[81]
  PIN crash_dump_o[80] 
    ANTENNAPARTIALMETALAREA 1.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.18 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 87.616 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.344 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 170.541 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[80]
  PIN crash_dump_o[79] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 34.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 128.168 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.9599 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 42.6646 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END crash_dump_o[79]
  PIN crash_dump_o[78] 
    ANTENNAPARTIALMETALAREA 1.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.292 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 46.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 174.048 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 41.4539 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 157.061 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.41844 LAYER VL ;
  END crash_dump_o[78]
  PIN crash_dump_o[77] 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 47.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 179.08 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.9855 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 60.6797 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER VL ;
  END crash_dump_o[77]
  PIN crash_dump_o[76] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 101.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 377.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.063 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 116.816 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02881 LAYER VL ;
  END crash_dump_o[76]
  PIN crash_dump_o[75] 
    ANTENNAPARTIALMETALAREA 0.84 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.256 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 54.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 201.872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.2421 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 68.9811 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[75]
  PIN crash_dump_o[74] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 62.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 233.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.3557 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 104.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER VL ;
  END crash_dump_o[74]
  PIN crash_dump_o[73] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 61.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 228.512 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.9703 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 75.3928 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02881 LAYER VL ;
  END crash_dump_o[73]
  PIN crash_dump_o[72] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 97.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 362.896 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.9357 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 105.266 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[72]
  PIN crash_dump_o[71] 
    ANTENNAPARTIALMETALAREA 2.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 97.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 364.672 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.1103 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 159.917 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER VL ;
  END crash_dump_o[71]
  PIN crash_dump_o[70] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 97.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 363.192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.8813 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 115.911 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END crash_dump_o[70]
  PIN crash_dump_o[69] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 59.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 220.52 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.0312 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 142.485 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER VL ;
  END crash_dump_o[69]
  PIN crash_dump_o[68] 
    ANTENNAPARTIALMETALAREA 0.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 86.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 322.344 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8656 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.51 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 102.897 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[68]
  PIN crash_dump_o[67] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 86.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 322.344 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8656 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.2693 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 90.9063 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[67]
  PIN crash_dump_o[66] 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 54.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 203.352 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8416 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.1685 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.273 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[66]
  PIN crash_dump_o[65] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 91.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 340.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8416 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.4334 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 113.18 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.806452 LAYER VL ;
  END crash_dump_o[65]
  PIN crash_dump_o[64] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 73.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 273.504 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8272 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.6603 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.5696 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER VL ;
  END crash_dump_o[64]
  PIN crash_dump_o[63] 
    ANTENNAPARTIALMETALAREA 0.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.96 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 44.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 165.168 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.88 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.7121 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 108.736 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[63]
  PIN crash_dump_o[62] 
    ANTENNAPARTIALMETALAREA 2.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 61.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 231.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.173 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 75.7896 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[62]
  PIN crash_dump_o[61] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 46.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 176.712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.4051 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 162.738 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[61]
  PIN crash_dump_o[60] 
    ANTENNAPARTIALMETALAREA 2.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 99.456 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.6473 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 78.0413 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[60]
  PIN crash_dump_o[59] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 70.744 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.3811 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 101.809 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[59]
  PIN crash_dump_o[58] 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 74.888 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.9969 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 61.7502 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[58]
  PIN crash_dump_o[57] 
    ANTENNAPARTIALMETALAREA 8.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.376 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 124.912 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.3992 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 66.5392 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[57]
  PIN crash_dump_o[56] 
    ANTENNAPARTIALMETALAREA 3.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.766 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 28.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 109.816 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.0267 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 77.43 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[56]
  PIN crash_dump_o[55] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.694 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 34.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 131.424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.5321 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 79.6305 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[55]
  PIN crash_dump_o[54] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.3262 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.064 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[54]
  PIN crash_dump_o[53] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 38.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 145.04 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.1351 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.936 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[53]
  PIN crash_dump_o[52] 
    ANTENNAPARTIALMETALAREA 1.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.292 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 49.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 189.44 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 43.9916 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 167.908 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[52]
  PIN crash_dump_o[51] 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 39 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 148.296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.1884 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 68.0344 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[51]
  PIN crash_dump_o[50] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 28.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 107.152 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.6999 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 117.902 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[50]
  PIN crash_dump_o[49] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 39.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 150.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.88 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.6955 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 172.072 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[49]
  PIN crash_dump_o[48] 
    ANTENNAPARTIALMETALAREA 0.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 100.936 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.8542 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 102.121 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[48]
  PIN crash_dump_o[47] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 51.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 195.656 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8344 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.5703 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 137.598 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.78571 LAYER VL ;
  END crash_dump_o[47]
  PIN crash_dump_o[46] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 33.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 128.168 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.9704 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 68.4212 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[46]
  PIN crash_dump_o[45] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 41.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 156.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8344 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.451 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 71.274 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.78571 LAYER VL ;
  END crash_dump_o[45]
  PIN crash_dump_o[44] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 42.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 159.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.591 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 105.58 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[44]
  PIN crash_dump_o[43] 
    ANTENNAPARTIALMETALAREA 3.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.838 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 60.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 229.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9616 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.3923 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 159.828 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[43]
  PIN crash_dump_o[42] 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.812 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 102.416 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.7816 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 60.1721 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[42]
  PIN crash_dump_o[41] 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 30.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 115.736 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.7574 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 82.3955 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[41]
  PIN crash_dump_o[40] 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.324 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 49.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 186.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.152 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 73.0185 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[40]
  PIN crash_dump_o[39] 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 38.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 145.928 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 56.2977 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 216.179 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END crash_dump_o[39]
  PIN crash_dump_o[38] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 49.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 186.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.1908 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 96.8497 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[38]
  PIN crash_dump_o[37] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 50.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 192.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9616 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.9655 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 138.679 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[37]
  PIN crash_dump_o[36] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 52.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 198.616 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.9325 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 153.107 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[36]
  PIN crash_dump_o[35] 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 56.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 208.976 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.88 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.1029 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 72.2845 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.41844 LAYER VL ;
  END crash_dump_o[35]
  PIN crash_dump_o[34] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 63.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 239.168 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.88 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.3395 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 123.393 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.41844 LAYER VL ;
  END crash_dump_o[34]
  PIN crash_dump_o[33] 
    ANTENNAPARTIALMETALAREA 0.92 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 58.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 217.264 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9712 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.2095 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 95.7402 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[33]
  PIN crash_dump_o[31] 
    ANTENNAPARTIALMETALAREA 0.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 96.792 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5872 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.5524 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 144.387 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.78571 LAYER VL ;
  END crash_dump_o[31]
  PIN crash_dump_o[30] 
    ANTENNAPARTIALMETALAREA 1.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.81 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 124.616 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5872 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.2485 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 121.311 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.78571 LAYER VL ;
  END crash_dump_o[30]
  PIN crash_dump_o[29] 
    ANTENNAPARTIALMETALAREA 1.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.928 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.8147 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 87.9154 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[29]
  PIN crash_dump_o[28] 
    ANTENNAPARTIALMETALAREA 5.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.312 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 120.01 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 445.785 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[28]
  PIN crash_dump_o[27] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 102.712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.3114 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 70.5572 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[27]
  PIN crash_dump_o[26] 
    ANTENNAPARTIALMETALAREA 21 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 77.996 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.304 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.8897 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 45.5396 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[26]
  PIN crash_dump_o[25] 
    ANTENNAPARTIALMETALAREA 2.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 97.088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.7824 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 72.4601 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[25]
  PIN crash_dump_o[24] 
    ANTENNAPARTIALMETALAREA 15.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 56.98 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.76187 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 37.6665 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[24]
  PIN crash_dump_o[23] 
    ANTENNAPARTIALMETALAREA 29.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 110.408 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.864 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.26394 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.5039 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[23]
  PIN crash_dump_o[22] 
    ANTENNAPARTIALMETALAREA 4.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.318 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.36 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.42513 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 33.0412 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[22]
  PIN crash_dump_o[21] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 30 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 113.96 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.2489 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 115.464 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[21]
  PIN crash_dump_o[20] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.68 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5872 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.6954 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 46.2252 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.78571 LAYER VL ;
  END crash_dump_o[20]
  PIN crash_dump_o[19] 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 82.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.87551 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 30.9275 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[19]
  PIN crash_dump_o[18] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 89.688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.6732 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 91.0118 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[18]
  PIN crash_dump_o[17] 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 34.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 131.128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.8372 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 45.7059 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[17]
  PIN crash_dump_o[16] 
    ANTENNAPARTIALMETALAREA 1.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.18 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 128.76 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.6747 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 45.0646 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[16]
  PIN crash_dump_o[15] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 33.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 126.392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5872 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.4411 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 157.187 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.38095 LAYER VL ;
  END crash_dump_o[15]
  PIN crash_dump_o[14] 
    ANTENNAPARTIALMETALAREA 1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.996 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 97.088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5872 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.292 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 58.4461 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.38095 LAYER VL ;
  END crash_dump_o[14]
  PIN crash_dump_o[13] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 37.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 140.6 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5872 LAYER M3 ; 
    ANTENNAMAXAREACAR 73.1544 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 283.897 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.7619 LAYER VL ;
  END crash_dump_o[13]
  PIN crash_dump_o[12] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 41.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 154.512 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.5304 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 138.39 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.62037 LAYER VL ;
  END crash_dump_o[12]
  PIN crash_dump_o[11] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 43.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 165.464 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.4242 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 51.578 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[11]
  PIN crash_dump_o[10] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 33.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 126.096 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5872 LAYER M3 ; 
    ANTENNAMAXAREACAR 72.7952 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 281.271 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.7619 LAYER VL ;
  END crash_dump_o[10]
  PIN crash_dump_o[9] 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 102.416 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5872 LAYER M3 ; 
    ANTENNAMAXAREACAR 62.4128 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 242.61 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VL ;
  END crash_dump_o[9]
  PIN crash_dump_o[8] 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 40.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 150.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.8798 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 49.2832 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[8]
  PIN crash_dump_o[7] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 35.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 134.976 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.6822 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 128.702 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END crash_dump_o[7]
  PIN crash_dump_o[6] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 46.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 174.048 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.5929 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 80.9488 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[6]
  PIN crash_dump_o[5] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 47.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 179.672 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.9487 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 57.1385 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[5]
  PIN crash_dump_o[4] 
    ANTENNAPARTIALMETALAREA 1.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.476 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 46.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 173.456 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.1671 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 145.14 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[4]
  PIN crash_dump_o[3] 
    ANTENNAPARTIALMETALAREA 0.84 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.256 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 39.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 148.592 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5872 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.6523 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 101.566 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.78571 LAYER VL ;
  END crash_dump_o[3]
  PIN crash_dump_o[2] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 43.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 163.984 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 56.9103 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 213.909 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[2]
  PIN crash_dump_o[1] 
    ANTENNAPARTIALMETALAREA 0.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 51.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 193.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.5118 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 154.699 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[1]
  PIN crash_dump_o[0] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 178.784 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.4936 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 92.8702 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[0]
  PIN double_fault_seen_o 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 41.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 155.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.9056 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.1026 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 67.4466 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0550661 LAYER VL ;
  END double_fault_seen_o
  PIN fetch_enable_i[3] 
  END fetch_enable_i[3]
  PIN fetch_enable_i[2] 
  END fetch_enable_i[2]
  PIN fetch_enable_i[1] 
  END fetch_enable_i[1]
  PIN fetch_enable_i[0] 
  END fetch_enable_i[0]
  PIN core_sleep_o 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 80.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 298.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.2066 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 104.59 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.606061 LAYER VL ;
  END core_sleep_o
  PIN scan_rst_ni 
  END scan_rst_ni
END ibex_top

END LIBRARY
