##
## LEF for PtnCells ;
## created by Innovus v19.10-p002_1 on Fri May 29 13:00:12 2020
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO mult8x8
  CLASS BLOCK ;
  SIZE 256.800000 BY 70.800000 ;
  FOREIGN mult8x8 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.14 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.666 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5544 LAYER M2  ;
    ANTENNAMAXAREACAR 20.5931 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 77.728 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER V2  ;
    ANTENNAMAXCUTCAR 1.22655 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 132.64 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 498.464 LAYER M3  ;
    ANTENNAGATEAREA 28.9728 LAYER M3  ;
    ANTENNAMAXAREACAR 25.1712 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 94.9325 LAYER M3  ;
    ANTENNAMAXCUTCAR 2.52525 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 11.900000 70.200000 12.100000 70.800000 ;
    END
  END clk
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.204 LAYER M2  ;
    ANTENNAMAXAREACAR 9.9451 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 36.9275 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.196078 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 23.900000 70.200000 24.100000 70.800000 ;
    END
  END resetn
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 26.7719 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 101.123 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 32.900000 0.600000 33.100000 ;
    END
  END a[7]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.06 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.622 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 28.9649 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 109.237 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 29.900000 0.600000 30.100000 ;
    END
  END a[6]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 24.1404 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 91.386 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 26.900000 0.600000 27.100000 ;
    END
  END a[5]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 30.2807 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 114.105 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 23.900000 0.600000 24.100000 ;
    END
  END a[4]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.26 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.362 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 27.6491 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 104.368 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 20.900000 0.600000 21.100000 ;
    END
  END a[3]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.98 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 24.5789 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 93.0088 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 17.900000 0.600000 18.100000 ;
    END
  END a[2]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.02 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.474 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 27.6491 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 104.368 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 14.900000 0.600000 15.100000 ;
    END
  END a[1]
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.06 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.622 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 27.2105 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 102.746 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 11.900000 0.600000 12.100000 ;
    END
  END a[0]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.42 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 29.4035 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 110.86 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 56.900000 0.600000 57.100000 ;
    END
  END b[7]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.14 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 26.3333 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 99.5 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 53.900000 0.600000 54.100000 ;
    END
  END b[6]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.26 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.362 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 31.1579 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 117.351 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 50.900000 0.600000 51.100000 ;
    END
  END b[5]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 25.4561 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 96.2544 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 47.900000 0.600000 48.100000 ;
    END
  END b[4]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.02 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.474 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3  ;
    ANTENNAMAXAREACAR 28.3468 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 107.189 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 44.900000 0.600000 45.100000 ;
    END
  END b[3]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 23.7018 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 89.7632 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 41.900000 0.600000 42.100000 ;
    END
  END b[2]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.586 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 23.2632 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 88.1404 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 38.900000 0.600000 39.100000 ;
    END
  END b[1]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.38 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.806 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 LAYER M3  ;
    ANTENNAMAXAREACAR 35.9825 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 135.202 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.31579 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 35.900000 0.600000 36.100000 ;
    END
  END b[0]
  PIN result[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.98 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.026 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.66 LAYER M3  ;
    ANTENNAMAXAREACAR 1.01389 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 3.80198 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.024024 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 56.900000 256.800000 57.100000 ;
    END
  END result[15]
  PIN result[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.62 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.242 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.603 LAYER M3  ;
    ANTENNAMAXAREACAR 2.07576 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 7.7841 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0461007 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 53.900000 256.800000 54.100000 ;
    END
  END result[14]
  PIN result[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.06 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.602 LAYER M3  ;
    ANTENNAMAXAREACAR 1.49716 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 5.63213 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0461184 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 50.900000 256.800000 51.100000 ;
    END
  END result[13]
  PIN result[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.47 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.603 LAYER M3  ;
    ANTENNAMAXAREACAR 1.58402 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 5.9078 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0461007 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 47.900000 256.800000 48.100000 ;
    END
  END result[12]
  PIN result[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.78 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.986 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.602 LAYER M3  ;
    ANTENNAMAXAREACAR 1.71238 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 6.42844 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0461184 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 44.900000 256.800000 45.100000 ;
    END
  END result[11]
  PIN result[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.02 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.174 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.603 LAYER M3  ;
    ANTENNAMAXAREACAR 1.46108 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 5.45294 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0461007 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 41.900000 256.800000 42.100000 ;
    END
  END result[10]
  PIN result[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.18 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.766 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.603 LAYER M3  ;
    ANTENNAMAXAREACAR 1.46108 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 5.45294 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0461007 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 38.900000 256.800000 39.100000 ;
    END
  END result[9]
  PIN result[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.99 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.602 LAYER M3  ;
    ANTENNAMAXAREACAR 1.29731 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 4.8927 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0461184 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 35.900000 256.800000 36.100000 ;
    END
  END result[8]
  PIN result[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.34 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.058 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.602 LAYER M3  ;
    ANTENNAMAXAREACAR 2.11207 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 7.9073 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0461184 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 32.900000 256.800000 33.100000 ;
    END
  END result[7]
  PIN result[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.34 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.358 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.893 LAYER M3  ;
    ANTENNAMAXAREACAR 2.21046 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 8.03212 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0845219 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 29.900000 256.800000 30.100000 ;
    END
  END result[6]
  PIN result[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.34 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.058 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.893 LAYER M3  ;
    ANTENNAMAXAREACAR 2.78098 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 10.1431 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0845219 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 26.900000 256.800000 27.100000 ;
    END
  END result[5]
  PIN result[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.18 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.466 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.848 LAYER M3  ;
    ANTENNAMAXAREACAR 1.94747 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 7.14466 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0561798 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 23.900000 256.800000 24.100000 ;
    END
  END result[4]
  PIN result[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.58 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.346 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.014 LAYER M3  ;
    ANTENNAMAXAREACAR 3.91976 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 14.6616 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0794439 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 20.900000 256.800000 21.100000 ;
    END
  END result[3]
  PIN result[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.78 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.386 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.014 LAYER M3  ;
    ANTENNAMAXAREACAR 3.6854 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 13.9168 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0794439 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 17.900000 256.800000 18.100000 ;
    END
  END result[2]
  PIN result[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.22 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.314 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.014 LAYER M3  ;
    ANTENNAMAXAREACAR 3.67349 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 14.03 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0794439 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 14.900000 256.800000 15.100000 ;
    END
  END result[1]
  PIN result[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.34 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.458 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.014 LAYER M3  ;
    ANTENNAMAXAREACAR 3.78073 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 14.1472 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0794439 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 256.200000 11.900000 256.800000 12.100000 ;
    END
  END result[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M3 ;
        RECT 1.200000 1.200000 255.600000 3.600000 ;
        RECT 1.200000 67.200000 255.600000 69.600000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M3 ;
        RECT 4.800000 4.800000 252.000000 7.200000 ;
        RECT 4.800000 63.600000 252.000000 66.000000 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 256.800000 70.800000 ;
    LAYER M2 ;
      RECT 26.020000 68.280000 256.800000 70.800000 ;
      RECT 14.020000 68.280000 21.980000 70.800000 ;
      RECT 0.000000 68.280000 9.980000 70.800000 ;
      RECT 0.000000 0.000000 256.800000 68.280000 ;
    LAYER M3 ;
      RECT 253.920000 61.680000 256.800000 65.280000 ;
      RECT 0.000000 61.680000 2.880000 65.280000 ;
      RECT 0.000000 59.020000 256.800000 61.680000 ;
      RECT 2.520000 9.980000 254.280000 59.020000 ;
      RECT 0.000000 9.120000 256.800000 9.980000 ;
      RECT 253.920000 5.520000 256.800000 9.120000 ;
      RECT 0.000000 5.520000 2.880000 9.120000 ;
  END
END mult8x8

END LIBRARY
