/homes/user/stud/fall23/yl5334/ibex_/ibex/mem_db/sram_top.lef