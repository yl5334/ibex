

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO ibex_top 
  PIN clk_i 
    ANTENNAPARTIALMETALAREA 3.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.578 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 43.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 161.912 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2352 LAYER M3 ; 
    ANTENNAMAXAREACAR 227.176 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 849.089 LAYER M3 ;
    ANTENNAMAXCUTCAR 5.55556 LAYER VL ;
  END clk_i
  PIN rst_ni 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END rst_ni
  PIN test_en_i 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.5721 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END test_en_i
  PIN ram_cfg_i[9] 
  END ram_cfg_i[9]
  PIN ram_cfg_i[8] 
  END ram_cfg_i[8]
  PIN ram_cfg_i[7] 
  END ram_cfg_i[7]
  PIN ram_cfg_i[6] 
  END ram_cfg_i[6]
  PIN ram_cfg_i[5] 
  END ram_cfg_i[5]
  PIN ram_cfg_i[4] 
  END ram_cfg_i[4]
  PIN ram_cfg_i[3] 
  END ram_cfg_i[3]
  PIN ram_cfg_i[2] 
  END ram_cfg_i[2]
  PIN ram_cfg_i[1] 
  END ram_cfg_i[1]
  PIN ram_cfg_i[0] 
  END ram_cfg_i[0]
  PIN hart_id_i[31] 
    ANTENNAPARTIALMETALAREA 3.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.482 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 146.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[31]
  PIN hart_id_i[30] 
    ANTENNAPARTIALMETALAREA 1.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.956 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.4189 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 98.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[30]
  PIN hart_id_i[29] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.806 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.6982 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 112.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[29]
  PIN hart_id_i[28] 
    ANTENNAPARTIALMETALAREA 2.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.844 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.9234 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[28]
  PIN hart_id_i[27] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.9324 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 57.1892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[27]
  PIN hart_id_i[26] 
    ANTENNAPARTIALMETALAREA 2.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.804 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.1306 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 141.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[26]
  PIN hart_id_i[25] 
    ANTENNAPARTIALMETALAREA 2.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.1757 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 123.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[25]
  PIN hart_id_i[24] 
    ANTENNAPARTIALMETALAREA 2.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.62 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.4279 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 131.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[24]
  PIN hart_id_i[23] 
    ANTENNAPARTIALMETALAREA 0.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.442 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.42793 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[23]
  PIN hart_id_i[22] 
    ANTENNAPARTIALMETALAREA 1.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.252 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.0225 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 111.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[22]
  PIN hart_id_i[21] 
    ANTENNAPARTIALMETALAREA 2.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.473 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 113.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[21]
  PIN hart_id_i[20] 
    ANTENNAPARTIALMETALAREA 2.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.436 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.1216 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 108.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[20]
  PIN hart_id_i[19] 
    ANTENNAPARTIALMETALAREA 2.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.7703 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[19]
  PIN hart_id_i[18] 
    ANTENNAPARTIALMETALAREA 1.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.956 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.518 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 94.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[18]
  PIN hart_id_i[17] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.9054 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 48.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[17]
  PIN hart_id_i[16] 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.0946 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 102.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[16]
  PIN hart_id_i[15] 
    ANTENNAPARTIALMETALAREA 2.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.5721 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[15]
  PIN hart_id_i[14] 
    ANTENNAPARTIALMETALAREA 2.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.028 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.9234 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[14]
  PIN hart_id_i[13] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.0676 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[13]
  PIN hart_id_i[12] 
    ANTENNAPARTIALMETALAREA 2.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.732 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.6261 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 124.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[12]
  PIN hart_id_i[11] 
    ANTENNAPARTIALMETALAREA 1.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.884 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.8604 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 68.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[11]
  PIN hart_id_i[10] 
    ANTENNAPARTIALMETALAREA 2.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.732 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.6261 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 124.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[10]
  PIN hart_id_i[9] 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.1757 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 123.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[9]
  PIN hart_id_i[8] 
    ANTENNAPARTIALMETALAREA 1.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.884 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.8604 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 68.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[8]
  PIN hart_id_i[7] 
    ANTENNAPARTIALMETALAREA 2.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.3739 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 116.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[7]
  PIN hart_id_i[6] 
    ANTENNAPARTIALMETALAREA 2.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.14 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.2207 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 104.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[6]
  PIN hart_id_i[5] 
    ANTENNAPARTIALMETALAREA 2.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.6712 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 106.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[5]
  PIN hart_id_i[4] 
    ANTENNAPARTIALMETALAREA 2.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.14 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.1216 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 108.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[4]
  PIN hart_id_i[3] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.545 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[3]
  PIN hart_id_i[2] 
    ANTENNAPARTIALMETALAREA 1.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.956 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.518 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 94.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[2]
  PIN hart_id_i[1] 
    ANTENNAPARTIALMETALAREA 2.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.6712 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 106.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[1]
  PIN hart_id_i[0] 
    ANTENNAPARTIALMETALAREA 1.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.956 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.0225 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 111.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END hart_id_i[0]
  PIN boot_addr_i[31] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.6441 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 98.8559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[31]
  PIN boot_addr_i[30] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[30]
  PIN boot_addr_i[29] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.8423 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 92.1892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[29]
  PIN boot_addr_i[28] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.622 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.4459 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 105.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[28]
  PIN boot_addr_i[27] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[27]
  PIN boot_addr_i[26] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.622 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.545 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 102.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[26]
  PIN boot_addr_i[25] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[25]
  PIN boot_addr_i[24] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.0676 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[24]
  PIN boot_addr_i[23] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.6712 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 106.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[23]
  PIN boot_addr_i[22] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[22]
  PIN boot_addr_i[21] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.622 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.545 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 102.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[21]
  PIN boot_addr_i[20] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[20]
  PIN boot_addr_i[19] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.545 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 102.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[19]
  PIN boot_addr_i[18] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.0676 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[18]
  PIN boot_addr_i[17] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[17]
  PIN boot_addr_i[16] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[16]
  PIN boot_addr_i[15] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[15]
  PIN boot_addr_i[14] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.6712 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 106.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[14]
  PIN boot_addr_i[13] 
    ANTENNAPARTIALMETALAREA 0.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.146 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.1667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 89.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[13]
  PIN boot_addr_i[12] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[12]
  PIN boot_addr_i[11] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.5225 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[11]
  PIN boot_addr_i[10] 
    ANTENNAPARTIALMETALAREA 0.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 8.97748 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 37.1892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END boot_addr_i[10]
  PIN boot_addr_i[9] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.2748 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 119.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[9]
  PIN boot_addr_i[8] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.8333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 153.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END boot_addr_i[8]
  PIN boot_addr_i[7] 
  END boot_addr_i[7]
  PIN boot_addr_i[6] 
  END boot_addr_i[6]
  PIN boot_addr_i[5] 
  END boot_addr_i[5]
  PIN boot_addr_i[4] 
  END boot_addr_i[4]
  PIN boot_addr_i[3] 
  END boot_addr_i[3]
  PIN boot_addr_i[2] 
  END boot_addr_i[2]
  PIN boot_addr_i[1] 
  END boot_addr_i[1]
  PIN boot_addr_i[0] 
  END boot_addr_i[0]
  PIN instr_req_o 
    ANTENNAPARTIALMETALAREA 7.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.676 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.7888 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.3396 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 70.2573 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.60417 LAYER VL ;
  END instr_req_o
  PIN instr_gnt_i 
    ANTENNAPARTIALMETALAREA 1.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.81 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.4369 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 73.8559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_gnt_i
  PIN instr_rvalid_i 
    ANTENNAPARTIALMETALAREA 0.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.182 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.5811 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 52.1892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rvalid_i
  PIN instr_addr_o[31] 
    ANTENNAPARTIALMETALAREA 1.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.736 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.965469 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.67156 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[31]
  PIN instr_addr_o[30] 
    ANTENNAPARTIALMETALAREA 2.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.508 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.35609 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.11687 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[30]
  PIN instr_addr_o[29] 
    ANTENNAPARTIALMETALAREA 0.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.37172 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.87469 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[29]
  PIN instr_addr_o[28] 
    ANTENNAPARTIALMETALAREA 7.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.084 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.05922 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 11.5919 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[28]
  PIN instr_addr_o[27] 
    ANTENNAPARTIALMETALAREA 1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.934219 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.55594 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[27]
  PIN instr_addr_o[26] 
    ANTENNAPARTIALMETALAREA 1.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.068 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.29359 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.88563 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[26]
  PIN instr_addr_o[25] 
    ANTENNAPARTIALMETALAREA 0.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.066 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.46266 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 16.7231 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.11257 LAYER VL ;
  END instr_addr_o[25]
  PIN instr_addr_o[24] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.066 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.84916 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 10.7531 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.150094 LAYER VL ;
  END instr_addr_o[24]
  PIN instr_addr_o[23] 
    ANTENNAPARTIALMETALAREA 1.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.066 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.21126 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.39287 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.11257 LAYER VL ;
  END instr_addr_o[23]
  PIN instr_addr_o[22] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.88734 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.0825 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[22]
  PIN instr_addr_o[21] 
    ANTENNAPARTIALMETALAREA 8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.896 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.69984 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.8466 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[21]
  PIN instr_addr_o[20] 
    ANTENNAPARTIALMETALAREA 7.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.564 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.12172 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 15.4075 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[20]
  PIN instr_addr_o[19] 
    ANTENNAPARTIALMETALAREA 0.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.934219 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.55594 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[19]
  PIN instr_addr_o[18] 
    ANTENNAPARTIALMETALAREA 0.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.13734 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.3075 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[18]
  PIN instr_addr_o[17] 
    ANTENNAPARTIALMETALAREA 0.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.066 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.46266 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 16.7231 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.11257 LAYER VL ;
  END instr_addr_o[17]
  PIN instr_addr_o[16] 
    ANTENNAPARTIALMETALAREA 0.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.404 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.606094 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2.34187 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[16]
  PIN instr_addr_o[15] 
    ANTENNAPARTIALMETALAREA 2.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.44984 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.52156 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[15]
  PIN instr_addr_o[14] 
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.48109 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.27937 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[14]
  PIN instr_addr_o[13] 
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.96 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.12172 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.24969 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[13]
  PIN instr_addr_o[12] 
    ANTENNAPARTIALMETALAREA 3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.692 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.21547 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.47 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[12]
  PIN instr_addr_o[11] 
    ANTENNAPARTIALMETALAREA 9.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.112 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.10609 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 15.3497 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[11]
  PIN instr_addr_o[10] 
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.88734 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.19813 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[10]
  PIN instr_addr_o[9] 
    ANTENNAPARTIALMETALAREA 0.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.15297 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.36531 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[9]
  PIN instr_addr_o[8] 
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.956 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.965469 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.72938 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[8]
  PIN instr_addr_o[7] 
    ANTENNAPARTIALMETALAREA 5.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.312 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.60609 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.79969 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[7]
  PIN instr_addr_o[6] 
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.01234 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 11.245 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[6]
  PIN instr_addr_o[5] 
    ANTENNAPARTIALMETALAREA 1.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.715469 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2.74656 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[5]
  PIN instr_addr_o[4] 
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.62 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.24672 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.77 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[4]
  PIN instr_addr_o[3] 
    ANTENNAPARTIALMETALAREA 2.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.90297 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 10.8403 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.046875 LAYER VL ;
  END instr_addr_o[3]
  PIN instr_addr_o[2] 
    ANTENNAPARTIALMETALAREA 0.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.746719 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2.92 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[2]
  PIN instr_rdata_i[31] 
    ANTENNAPARTIALMETALAREA 1.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.402 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.8423 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.8559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[31]
  PIN instr_rdata_i[30] 
    ANTENNAPARTIALMETALAREA 0.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.4009 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 125.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[30]
  PIN instr_rdata_i[29] 
    ANTENNAPARTIALMETALAREA 1.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.106 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.9414 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 90.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[29]
  PIN instr_rdata_i[28] 
    ANTENNAPARTIALMETALAREA 0.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.294 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.5541 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 135.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[28]
  PIN instr_rdata_i[27] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.474 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.1486 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 117.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[27]
  PIN instr_rdata_i[26] 
    ANTENNAPARTIALMETALAREA 0.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.6982 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 115.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[26]
  PIN instr_rdata_i[25] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.8964 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 107.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[25]
  PIN instr_rdata_i[24] 
    ANTENNAPARTIALMETALAREA 0.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.527 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 126.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[24]
  PIN instr_rdata_i[23] 
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.146 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.2027 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 130.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[23]
  PIN instr_rdata_i[22] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.0495 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 118.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[22]
  PIN instr_rdata_i[21] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.258 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.7973 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[21]
  PIN instr_rdata_i[20] 
    ANTENNAPARTIALMETALAREA 0.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.2477 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 112.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[20]
  PIN instr_rdata_i[19] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.258 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.5991 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 117.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[19]
  PIN instr_rdata_i[18] 
    ANTENNAPARTIALMETALAREA 0.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.886 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.7793 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 45.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[18]
  PIN instr_rdata_i[17] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.8964 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 107.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[17]
  PIN instr_rdata_i[16] 
    ANTENNAPARTIALMETALAREA 0.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.9505 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 122.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[16]
  PIN instr_rdata_i[15] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.7973 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[15]
  PIN instr_rdata_i[14] 
    ANTENNAPARTIALMETALAREA 0.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.1486 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 115.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[14]
  PIN instr_rdata_i[13] 
    ANTENNAPARTIALMETALAREA 0.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.442 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.7523 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 130.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[13]
  PIN instr_rdata_i[12] 
    ANTENNAPARTIALMETALAREA 0.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.406 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.2477 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 112.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[12]
  PIN instr_rdata_i[11] 
    ANTENNAPARTIALMETALAREA 0.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.442 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.6532 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 133.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[11]
  PIN instr_rdata_i[10] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.622 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.6441 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 102.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[10]
  PIN instr_rdata_i[9] 
    ANTENNAPARTIALMETALAREA 0.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.554 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.6982 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 113.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[9]
  PIN instr_rdata_i[8] 
    ANTENNAPARTIALMETALAREA 0.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.1486 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 115.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[8]
  PIN instr_rdata_i[7] 
    ANTENNAPARTIALMETALAREA 0.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.554 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.0495 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 120.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[7]
  PIN instr_rdata_i[6] 
    ANTENNAPARTIALMETALAREA 1.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.366 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.6892 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 82.1892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[6]
  PIN instr_rdata_i[5] 
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.146 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.4009 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 123.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[5]
  PIN instr_rdata_i[4] 
    ANTENNAPARTIALMETALAREA 1.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.366 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.6892 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 82.1892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[4]
  PIN instr_rdata_i[3] 
    ANTENNAPARTIALMETALAREA 1.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.514 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.6351 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 67.1892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[3]
  PIN instr_rdata_i[2] 
    ANTENNAPARTIALMETALAREA 0.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.5721 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_rdata_i[2]
  PIN instr_rdata_i[1] 
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.6441 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 100.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[1]
  PIN instr_rdata_i[0] 
    ANTENNAPARTIALMETALAREA 0.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.294 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.5541 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 135.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_rdata_i[0]
  PIN instr_rdata_intg_i[6] 
  END instr_rdata_intg_i[6]
  PIN instr_rdata_intg_i[5] 
  END instr_rdata_intg_i[5]
  PIN instr_rdata_intg_i[4] 
  END instr_rdata_intg_i[4]
  PIN instr_rdata_intg_i[3] 
  END instr_rdata_intg_i[3]
  PIN instr_rdata_intg_i[2] 
  END instr_rdata_intg_i[2]
  PIN instr_rdata_intg_i[1] 
  END instr_rdata_intg_i[1]
  PIN instr_rdata_intg_i[0] 
  END instr_rdata_intg_i[0]
  PIN instr_err_i 
    ANTENNAPARTIALMETALAREA 1.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.662 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.7883 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 78.8559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END instr_err_i
  PIN data_req_o 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.252 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.944 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.488 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.47926 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.48842 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0482315 LAYER VL ;
  END data_req_o
  PIN data_gnt_i 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.95045 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 29.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_gnt_i
  PIN data_rvalid_i 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.95045 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 29.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rvalid_i
  PIN data_we_o 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 114.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 425.352 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2796 LAYER M3 ; 
    ANTENNAMAXAREACAR 41.5456 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 157.807 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END data_we_o
  PIN data_be_o[3] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.16 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.90414 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 25.5734 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.137931 LAYER VL ;
  END data_be_o[3]
  PIN data_be_o[2] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.862 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.06842 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.67666 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0197824 LAYER VL ;
  END data_be_o[2]
  PIN data_be_o[1] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.066 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.77373 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 15.3887 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0750469 LAYER V2 ;
  END data_be_o[1]
  PIN data_be_o[0] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.182 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.046 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.704008 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2.77146 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.058651 LAYER VL ;
  END data_be_o[0]
  PIN data_addr_o[31] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 83.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8464 LAYER M3 ; 
    ANTENNAMAXAREACAR 91.8817 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 356.231 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.78571 LAYER VL ;
  END data_addr_o[31]
  PIN data_addr_o[30] 
    ANTENNAPARTIALMETALAREA 1.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.512 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 61.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 231.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3664 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.3256 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 155.572 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.87356 LAYER VL ;
  END data_addr_o[30]
  PIN data_addr_o[29] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 65.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 244.792 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4164 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.6934 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 126.012 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.93798 LAYER VL ;
  END data_addr_o[29]
  PIN data_addr_o[28] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 73.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 275.872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4884 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.3437 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 136.311 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.16279 LAYER VL ;
  END data_addr_o[28]
  PIN data_addr_o[27] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 69.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 258.704 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9088 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.2655 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 85.1496 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.41844 LAYER VL ;
  END data_addr_o[27]
  PIN data_addr_o[26] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 54.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 205.424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9088 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.773 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 104.046 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.16279 LAYER VL ;
  END data_addr_o[26]
  PIN data_addr_o[25] 
    ANTENNAPARTIALMETALAREA 1.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.18 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 64.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 239.168 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9088 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.7001 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 100.78 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.16279 LAYER VL ;
  END data_addr_o[25]
  PIN data_addr_o[24] 
    ANTENNAPARTIALMETALAREA 2.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 87.912 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3664 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.6343 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 55.6875 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.72414 LAYER VL ;
  END data_addr_o[24]
  PIN data_addr_o[23] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 156.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9088 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.5893 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 66.024 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.16279 LAYER VL ;
  END data_addr_o[23]
  PIN data_addr_o[22] 
    ANTENNAPARTIALMETALAREA 0.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 59.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 223.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4164 LAYER M3 ; 
    ANTENNAMAXAREACAR 94.8941 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 365.886 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END data_addr_o[22]
  PIN data_addr_o[21] 
    ANTENNAPARTIALMETALAREA 4.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.428 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 90 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 335.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9664 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.6906 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 179.544 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END data_addr_o[21]
  PIN data_addr_o[20] 
    ANTENNAPARTIALMETALAREA 1.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.736 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 67.488 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1936 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.6071 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 53.684 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.87356 LAYER VL ;
  END data_addr_o[20]
  PIN data_addr_o[19] 
    ANTENNAPARTIALMETALAREA 1.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.144 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 69.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 258.852 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9088 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.6629 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.374 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.16279 LAYER VL ;
  END data_addr_o[19]
  PIN data_addr_o[18] 
    ANTENNAPARTIALMETALAREA 0.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 41.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 155.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3664 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.0229 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 136.263 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.23478 LAYER VL ;
  END data_addr_o[18]
  PIN data_addr_o[17] 
    ANTENNAPARTIALMETALAREA 1.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.66 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 61.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 231.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4164 LAYER M3 ; 
    ANTENNAMAXAREACAR 41.3625 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 158.784 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END data_addr_o[17]
  PIN data_addr_o[16] 
    ANTENNAPARTIALMETALAREA 1.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.736 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 89.688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3664 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.1379 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 198.57 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END data_addr_o[16]
  PIN data_addr_o[15] 
    ANTENNAPARTIALMETALAREA 0.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 40.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 150.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3664 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.9568 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 64.2668 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.16279 LAYER VL ;
  END data_addr_o[15]
  PIN data_addr_o[14] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 43.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 164.576 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5392 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.6595 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 90.1691 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.16279 LAYER VL ;
  END data_addr_o[14]
  PIN data_addr_o[13] 
    ANTENNAPARTIALMETALAREA 1.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.66 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 61.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 228.216 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2368 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.0901 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 143.255 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.77305 LAYER VL ;
  END data_addr_o[13]
  PIN data_addr_o[12] 
    ANTENNAPARTIALMETALAREA 1.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.144 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 38.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 142.08 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2368 LAYER M3 ; 
    ANTENNAMAXAREACAR 48.0336 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 178.566 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.55039 LAYER VL ;
  END data_addr_o[12]
  PIN data_addr_o[11] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 104.192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1936 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.6659 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 43.9625 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.16279 LAYER VL ;
  END data_addr_o[11]
  PIN data_addr_o[10] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 98.568 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3064 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.7248 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 117.352 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.87356 LAYER VL ;
  END data_addr_o[10]
  PIN data_addr_o[9] 
    ANTENNAPARTIALMETALAREA 2.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.396 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 52.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 199.8 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2584 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.9394 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 75.5239 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.16279 LAYER VL ;
  END data_addr_o[9]
  PIN data_addr_o[8] 
    ANTENNAPARTIALMETALAREA 2.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 122.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.1129 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 145.341 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.12766 LAYER VL ;
  END data_addr_o[8]
  PIN data_addr_o[7] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 100.048 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2128 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.4947 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 115.589 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.93798 LAYER VL ;
  END data_addr_o[7]
  PIN data_addr_o[6] 
    ANTENNAPARTIALMETALAREA 0.92 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 34.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 129.056 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3856 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.6488 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 99.2705 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END data_addr_o[6]
  PIN data_addr_o[5] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 44.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 167.536 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8488 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.6523 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 75.3166 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.16279 LAYER VL ;
  END data_addr_o[5]
  PIN data_addr_o[4] 
    ANTENNAPARTIALMETALAREA 1.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.92 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 61.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 230.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9304 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.9295 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 78.5334 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.16279 LAYER VL ;
  END data_addr_o[4]
  PIN data_addr_o[3] 
    ANTENNAPARTIALMETALAREA 2.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.028 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 31.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 120.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3856 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.4488 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 98.558 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.15054 LAYER VL ;
  END data_addr_o[3]
  PIN data_addr_o[2] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 74.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 279.128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9304 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.6459 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 85.2231 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.16279 LAYER VL ;
  END data_addr_o[2]
  PIN data_wdata_o[31] 
    ANTENNAPARTIALMETALAREA 1.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.292 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.95303 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.44583 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[31]
  PIN data_wdata_o[30] 
    ANTENNAPARTIALMETALAREA 0.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.50417 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 6.02822 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER V2 ;
  END data_wdata_o[30]
  PIN data_wdata_o[29] 
    ANTENNAPARTIALMETALAREA 1.68 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.364 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.864 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.44167 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 16.9875 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[29]
  PIN data_wdata_o[28] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.19545 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 23.4799 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[28]
  PIN data_wdata_o[27] 
    ANTENNAPARTIALMETALAREA 0.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.152 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.23712 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 20.2678 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[27]
  PIN data_wdata_o[26] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.728 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.96742 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.42424 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[26]
  PIN data_wdata_o[25] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 56.24 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.32727 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 27.7462 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[25]
  PIN data_wdata_o[24] 
    ANTENNAPARTIALMETALAREA 1.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.144 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.6303 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.94697 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[24]
  PIN data_wdata_o[23] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.38864 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 5.58409 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER V2 ;
  END data_wdata_o[23]
  PIN data_wdata_o[22] 
    ANTENNAPARTIALMETALAREA 1.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.624 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.09621 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.20076 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[22]
  PIN data_wdata_o[21] 
    ANTENNAPARTIALMETALAREA 1.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.66 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.28 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.03258 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 11.5102 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[21]
  PIN data_wdata_o[20] 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.64242 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 21.5405 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[20]
  PIN data_wdata_o[19] 
    ANTENNAPARTIALMETALAREA 2.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.916 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.976 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.86212 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 14.8966 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[19]
  PIN data_wdata_o[18] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.64 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.29318 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 31.25 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[18]
  PIN data_wdata_o[17] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.504 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.79697 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 25.6439 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[17]
  PIN data_wdata_o[16] 
    ANTENNAPARTIALMETALAREA 0.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.01364 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.53674 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[16]
  PIN data_wdata_o[15] 
    ANTENNAPARTIALMETALAREA 1.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.884 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.25606 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 4.8303 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER V2 ;
  END data_wdata_o[15]
  PIN data_wdata_o[14] 
    ANTENNAPARTIALMETALAREA 1.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.328 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.68 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.52045 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.3106 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[14]
  PIN data_wdata_o[13] 
    ANTENNAPARTIALMETALAREA 1.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.656 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.00606 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.52538 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[13]
  PIN data_wdata_o[12] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.224 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.01742 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 18.7489 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[12]
  PIN data_wdata_o[11] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.32 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.42197 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.10606 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[11]
  PIN data_wdata_o[10] 
    ANTENNAPARTIALMETALAREA 1.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.92 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.52 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.07045 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 19.1239 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[10]
  PIN data_wdata_o[9] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.208 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.47879 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.38636 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[9]
  PIN data_wdata_o[8] 
    ANTENNAPARTIALMETALAREA 0.92 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.552 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.025 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.94205 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER V2 ;
  END data_wdata_o[8]
  PIN data_wdata_o[7] 
    ANTENNAPARTIALMETALAREA 1.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.66 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.504 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.68788 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 10.4117 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[7]
  PIN data_wdata_o[6] 
    ANTENNAPARTIALMETALAREA 2.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.344 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.57727 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.7311 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[6]
  PIN data_wdata_o[5] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.976 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.09697 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 15.5784 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[5]
  PIN data_wdata_o[4] 
    ANTENNAPARTIALMETALAREA 2.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.34242 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 5.04167 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0189394 LAYER V2 ;
  END data_wdata_o[4]
  PIN data_wdata_o[3] 
    ANTENNAPARTIALMETALAREA 2.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.028 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.584848 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2.23864 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0568182 LAYER VL ;
  END data_wdata_o[3]
  PIN data_wdata_o[2] 
    ANTENNAPARTIALMETALAREA 0.68 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.6803 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.9269 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[2]
  PIN data_wdata_o[1] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.85758 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 11.2902 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[1]
  PIN data_wdata_o[0] 
    ANTENNAPARTIALMETALAREA 1.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.736 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.45303 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.58598 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0757576 LAYER VL ;
  END data_wdata_o[0]
  PIN data_rdata_i[31] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.7432 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 95.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[31]
  PIN data_rdata_i[30] 
    ANTENNAPARTIALMETALAREA 0.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 6.72523 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 28.8559 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[30]
  PIN data_rdata_i[29] 
    ANTENNAPARTIALMETALAREA 0.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.146 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.9775 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 129.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[29]
  PIN data_rdata_i[28] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.7432 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 95.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[28]
  PIN data_rdata_i[27] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.5721 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[27]
  PIN data_rdata_i[26] 
    ANTENNAPARTIALMETALAREA 0.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 6.72523 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 28.8559 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[26]
  PIN data_rdata_i[25] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 41.1847 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 156.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[25]
  PIN data_rdata_i[24] 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.8784 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 133.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[24]
  PIN data_rdata_i[23] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.2838 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 153.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[23]
  PIN data_rdata_i[22] 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.6441 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 98.8559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[22]
  PIN data_rdata_i[21] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.2748 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 119.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[21]
  PIN data_rdata_i[20] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.7432 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 95.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[20]
  PIN data_rdata_i[19] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.656 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.5811 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 143.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[19]
  PIN data_rdata_i[18] 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.806 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.1486 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 115.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[18]
  PIN data_rdata_i[17] 
    ANTENNAPARTIALMETALAREA 0.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 8.97748 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 37.1892 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[17]
  PIN data_rdata_i[16] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.473 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 113.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[16]
  PIN data_rdata_i[15] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.7703 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[15]
  PIN data_rdata_i[14] 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.482 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 146.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[14]
  PIN data_rdata_i[13] 
    ANTENNAPARTIALMETALAREA 1.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.476 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.3559 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 49.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[13]
  PIN data_rdata_i[12] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.8333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 153.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[12]
  PIN data_rdata_i[11] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.7432 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 95.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[11]
  PIN data_rdata_i[10] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.544 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.0315 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 146.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[10]
  PIN data_rdata_i[9] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.4459 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 105.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[9]
  PIN data_rdata_i[8] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.7432 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 95.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[8]
  PIN data_rdata_i[7] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.8423 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 92.1892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[7]
  PIN data_rdata_i[6] 
    ANTENNAPARTIALMETALAREA 0.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 6.72523 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 28.8559 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END data_rdata_i[6]
  PIN data_rdata_i[5] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.8423 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 92.1892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[5]
  PIN data_rdata_i[4] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.3739 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 116.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[4]
  PIN data_rdata_i[3] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.5721 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[3]
  PIN data_rdata_i[2] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.95045 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 29.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[2]
  PIN data_rdata_i[1] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.8423 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 92.1892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[1]
  PIN data_rdata_i[0] 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.9685 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 96.3559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_rdata_i[0]
  PIN data_rdata_intg_i[6] 
  END data_rdata_intg_i[6]
  PIN data_rdata_intg_i[5] 
  END data_rdata_intg_i[5]
  PIN data_rdata_intg_i[4] 
  END data_rdata_intg_i[4]
  PIN data_rdata_intg_i[3] 
  END data_rdata_intg_i[3]
  PIN data_rdata_intg_i[2] 
  END data_rdata_intg_i[2]
  PIN data_rdata_intg_i[1] 
  END data_rdata_intg_i[1]
  PIN data_rdata_intg_i[0] 
  END data_rdata_intg_i[0]
  PIN data_err_i 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.8423 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 92.1892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END data_err_i
  PIN irq_software_i 
    ANTENNAPARTIALMETALAREA 1.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.586 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.8423 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 90.5225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_software_i
  PIN irq_timer_i 
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.1667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 89.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_timer_i
  PIN irq_external_i 
    ANTENNAPARTIALMETALAREA 2.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.916 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.0766 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 128.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_external_i
  PIN irq_fast_i[14] 
    ANTENNAPARTIALMETALAREA 2.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.916 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.3288 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 134.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[14]
  PIN irq_fast_i[13] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.3559 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 140.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[13]
  PIN irq_fast_i[12] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.7342 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 63.8559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[12]
  PIN irq_fast_i[11] 
    ANTENNAPARTIALMETALAREA 2.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.844 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.527 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 128.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[11]
  PIN irq_fast_i[10] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.8063 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 51.3559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[10]
  PIN irq_fast_i[9] 
    ANTENNAPARTIALMETALAREA 2.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.732 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.4279 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 131.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[9]
  PIN irq_fast_i[8] 
    ANTENNAPARTIALMETALAREA 2.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.804 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.3288 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 134.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[8]
  PIN irq_fast_i[7] 
    ANTENNAPARTIALMETALAREA 2.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.73 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.3649 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 173.856 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[7]
  PIN irq_fast_i[6] 
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.7793 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 136.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[6]
  PIN irq_fast_i[5] 
    ANTENNAPARTIALMETALAREA 1.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.956 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.4189 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 98.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[5]
  PIN irq_fast_i[4] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.9685 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 96.3559 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[4]
  PIN irq_fast_i[3] 
    ANTENNAPARTIALMETALAREA 1.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.586 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.3468 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 107.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[3]
  PIN irq_fast_i[2] 
    ANTENNAPARTIALMETALAREA 1.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.8694 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 99.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[2]
  PIN irq_fast_i[1] 
    ANTENNAPARTIALMETALAREA 2.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.324 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.8243 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 118.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[1]
  PIN irq_fast_i[0] 
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.1667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 89.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_fast_i[0]
  PIN irq_nm_i 
    ANTENNAPARTIALMETALAREA 2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.548 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.2207 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 104.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END irq_nm_i
  PIN scramble_key_valid_i 
  END scramble_key_valid_i
  PIN scramble_key_i[127] 
  END scramble_key_i[127]
  PIN scramble_key_i[126] 
  END scramble_key_i[126]
  PIN scramble_key_i[125] 
  END scramble_key_i[125]
  PIN scramble_key_i[124] 
  END scramble_key_i[124]
  PIN scramble_key_i[123] 
  END scramble_key_i[123]
  PIN scramble_key_i[122] 
  END scramble_key_i[122]
  PIN scramble_key_i[121] 
  END scramble_key_i[121]
  PIN scramble_key_i[120] 
  END scramble_key_i[120]
  PIN scramble_key_i[119] 
  END scramble_key_i[119]
  PIN scramble_key_i[118] 
  END scramble_key_i[118]
  PIN scramble_key_i[117] 
  END scramble_key_i[117]
  PIN scramble_key_i[116] 
  END scramble_key_i[116]
  PIN scramble_key_i[115] 
  END scramble_key_i[115]
  PIN scramble_key_i[114] 
  END scramble_key_i[114]
  PIN scramble_key_i[113] 
  END scramble_key_i[113]
  PIN scramble_key_i[112] 
  END scramble_key_i[112]
  PIN scramble_key_i[111] 
  END scramble_key_i[111]
  PIN scramble_key_i[110] 
  END scramble_key_i[110]
  PIN scramble_key_i[109] 
  END scramble_key_i[109]
  PIN scramble_key_i[108] 
  END scramble_key_i[108]
  PIN scramble_key_i[107] 
  END scramble_key_i[107]
  PIN scramble_key_i[106] 
  END scramble_key_i[106]
  PIN scramble_key_i[105] 
  END scramble_key_i[105]
  PIN scramble_key_i[104] 
  END scramble_key_i[104]
  PIN scramble_key_i[103] 
  END scramble_key_i[103]
  PIN scramble_key_i[102] 
  END scramble_key_i[102]
  PIN scramble_key_i[101] 
  END scramble_key_i[101]
  PIN scramble_key_i[100] 
  END scramble_key_i[100]
  PIN scramble_key_i[99] 
  END scramble_key_i[99]
  PIN scramble_key_i[98] 
  END scramble_key_i[98]
  PIN scramble_key_i[97] 
  END scramble_key_i[97]
  PIN scramble_key_i[96] 
  END scramble_key_i[96]
  PIN scramble_key_i[95] 
  END scramble_key_i[95]
  PIN scramble_key_i[94] 
  END scramble_key_i[94]
  PIN scramble_key_i[93] 
  END scramble_key_i[93]
  PIN scramble_key_i[92] 
  END scramble_key_i[92]
  PIN scramble_key_i[91] 
  END scramble_key_i[91]
  PIN scramble_key_i[90] 
  END scramble_key_i[90]
  PIN scramble_key_i[89] 
  END scramble_key_i[89]
  PIN scramble_key_i[88] 
  END scramble_key_i[88]
  PIN scramble_key_i[87] 
  END scramble_key_i[87]
  PIN scramble_key_i[86] 
  END scramble_key_i[86]
  PIN scramble_key_i[85] 
  END scramble_key_i[85]
  PIN scramble_key_i[84] 
  END scramble_key_i[84]
  PIN scramble_key_i[83] 
  END scramble_key_i[83]
  PIN scramble_key_i[82] 
  END scramble_key_i[82]
  PIN scramble_key_i[81] 
  END scramble_key_i[81]
  PIN scramble_key_i[80] 
  END scramble_key_i[80]
  PIN scramble_key_i[79] 
  END scramble_key_i[79]
  PIN scramble_key_i[78] 
  END scramble_key_i[78]
  PIN scramble_key_i[77] 
  END scramble_key_i[77]
  PIN scramble_key_i[76] 
  END scramble_key_i[76]
  PIN scramble_key_i[75] 
  END scramble_key_i[75]
  PIN scramble_key_i[74] 
  END scramble_key_i[74]
  PIN scramble_key_i[73] 
  END scramble_key_i[73]
  PIN scramble_key_i[72] 
  END scramble_key_i[72]
  PIN scramble_key_i[71] 
  END scramble_key_i[71]
  PIN scramble_key_i[70] 
  END scramble_key_i[70]
  PIN scramble_key_i[69] 
  END scramble_key_i[69]
  PIN scramble_key_i[68] 
  END scramble_key_i[68]
  PIN scramble_key_i[67] 
  END scramble_key_i[67]
  PIN scramble_key_i[66] 
  END scramble_key_i[66]
  PIN scramble_key_i[65] 
  END scramble_key_i[65]
  PIN scramble_key_i[64] 
  END scramble_key_i[64]
  PIN scramble_key_i[63] 
  END scramble_key_i[63]
  PIN scramble_key_i[62] 
  END scramble_key_i[62]
  PIN scramble_key_i[61] 
  END scramble_key_i[61]
  PIN scramble_key_i[60] 
  END scramble_key_i[60]
  PIN scramble_key_i[59] 
  END scramble_key_i[59]
  PIN scramble_key_i[58] 
  END scramble_key_i[58]
  PIN scramble_key_i[57] 
  END scramble_key_i[57]
  PIN scramble_key_i[56] 
  END scramble_key_i[56]
  PIN scramble_key_i[55] 
  END scramble_key_i[55]
  PIN scramble_key_i[54] 
  END scramble_key_i[54]
  PIN scramble_key_i[53] 
  END scramble_key_i[53]
  PIN scramble_key_i[52] 
  END scramble_key_i[52]
  PIN scramble_key_i[51] 
  END scramble_key_i[51]
  PIN scramble_key_i[50] 
  END scramble_key_i[50]
  PIN scramble_key_i[49] 
  END scramble_key_i[49]
  PIN scramble_key_i[48] 
  END scramble_key_i[48]
  PIN scramble_key_i[47] 
  END scramble_key_i[47]
  PIN scramble_key_i[46] 
  END scramble_key_i[46]
  PIN scramble_key_i[45] 
  END scramble_key_i[45]
  PIN scramble_key_i[44] 
  END scramble_key_i[44]
  PIN scramble_key_i[43] 
  END scramble_key_i[43]
  PIN scramble_key_i[42] 
  END scramble_key_i[42]
  PIN scramble_key_i[41] 
  END scramble_key_i[41]
  PIN scramble_key_i[40] 
  END scramble_key_i[40]
  PIN scramble_key_i[39] 
  END scramble_key_i[39]
  PIN scramble_key_i[38] 
  END scramble_key_i[38]
  PIN scramble_key_i[37] 
  END scramble_key_i[37]
  PIN scramble_key_i[36] 
  END scramble_key_i[36]
  PIN scramble_key_i[35] 
  END scramble_key_i[35]
  PIN scramble_key_i[34] 
  END scramble_key_i[34]
  PIN scramble_key_i[33] 
  END scramble_key_i[33]
  PIN scramble_key_i[32] 
  END scramble_key_i[32]
  PIN scramble_key_i[31] 
  END scramble_key_i[31]
  PIN scramble_key_i[30] 
  END scramble_key_i[30]
  PIN scramble_key_i[29] 
  END scramble_key_i[29]
  PIN scramble_key_i[28] 
  END scramble_key_i[28]
  PIN scramble_key_i[27] 
  END scramble_key_i[27]
  PIN scramble_key_i[26] 
  END scramble_key_i[26]
  PIN scramble_key_i[25] 
  END scramble_key_i[25]
  PIN scramble_key_i[24] 
  END scramble_key_i[24]
  PIN scramble_key_i[23] 
  END scramble_key_i[23]
  PIN scramble_key_i[22] 
  END scramble_key_i[22]
  PIN scramble_key_i[21] 
  END scramble_key_i[21]
  PIN scramble_key_i[20] 
  END scramble_key_i[20]
  PIN scramble_key_i[19] 
  END scramble_key_i[19]
  PIN scramble_key_i[18] 
  END scramble_key_i[18]
  PIN scramble_key_i[17] 
  END scramble_key_i[17]
  PIN scramble_key_i[16] 
  END scramble_key_i[16]
  PIN scramble_key_i[15] 
  END scramble_key_i[15]
  PIN scramble_key_i[14] 
  END scramble_key_i[14]
  PIN scramble_key_i[13] 
  END scramble_key_i[13]
  PIN scramble_key_i[12] 
  END scramble_key_i[12]
  PIN scramble_key_i[11] 
  END scramble_key_i[11]
  PIN scramble_key_i[10] 
  END scramble_key_i[10]
  PIN scramble_key_i[9] 
  END scramble_key_i[9]
  PIN scramble_key_i[8] 
  END scramble_key_i[8]
  PIN scramble_key_i[7] 
  END scramble_key_i[7]
  PIN scramble_key_i[6] 
  END scramble_key_i[6]
  PIN scramble_key_i[5] 
  END scramble_key_i[5]
  PIN scramble_key_i[4] 
  END scramble_key_i[4]
  PIN scramble_key_i[3] 
  END scramble_key_i[3]
  PIN scramble_key_i[2] 
  END scramble_key_i[2]
  PIN scramble_key_i[1] 
  END scramble_key_i[1]
  PIN scramble_key_i[0] 
  END scramble_key_i[0]
  PIN scramble_nonce_i[63] 
  END scramble_nonce_i[63]
  PIN scramble_nonce_i[62] 
  END scramble_nonce_i[62]
  PIN scramble_nonce_i[61] 
  END scramble_nonce_i[61]
  PIN scramble_nonce_i[60] 
  END scramble_nonce_i[60]
  PIN scramble_nonce_i[59] 
  END scramble_nonce_i[59]
  PIN scramble_nonce_i[58] 
  END scramble_nonce_i[58]
  PIN scramble_nonce_i[57] 
  END scramble_nonce_i[57]
  PIN scramble_nonce_i[56] 
  END scramble_nonce_i[56]
  PIN scramble_nonce_i[55] 
  END scramble_nonce_i[55]
  PIN scramble_nonce_i[54] 
  END scramble_nonce_i[54]
  PIN scramble_nonce_i[53] 
  END scramble_nonce_i[53]
  PIN scramble_nonce_i[52] 
  END scramble_nonce_i[52]
  PIN scramble_nonce_i[51] 
  END scramble_nonce_i[51]
  PIN scramble_nonce_i[50] 
  END scramble_nonce_i[50]
  PIN scramble_nonce_i[49] 
  END scramble_nonce_i[49]
  PIN scramble_nonce_i[48] 
  END scramble_nonce_i[48]
  PIN scramble_nonce_i[47] 
  END scramble_nonce_i[47]
  PIN scramble_nonce_i[46] 
  END scramble_nonce_i[46]
  PIN scramble_nonce_i[45] 
  END scramble_nonce_i[45]
  PIN scramble_nonce_i[44] 
  END scramble_nonce_i[44]
  PIN scramble_nonce_i[43] 
  END scramble_nonce_i[43]
  PIN scramble_nonce_i[42] 
  END scramble_nonce_i[42]
  PIN scramble_nonce_i[41] 
  END scramble_nonce_i[41]
  PIN scramble_nonce_i[40] 
  END scramble_nonce_i[40]
  PIN scramble_nonce_i[39] 
  END scramble_nonce_i[39]
  PIN scramble_nonce_i[38] 
  END scramble_nonce_i[38]
  PIN scramble_nonce_i[37] 
  END scramble_nonce_i[37]
  PIN scramble_nonce_i[36] 
  END scramble_nonce_i[36]
  PIN scramble_nonce_i[35] 
  END scramble_nonce_i[35]
  PIN scramble_nonce_i[34] 
  END scramble_nonce_i[34]
  PIN scramble_nonce_i[33] 
  END scramble_nonce_i[33]
  PIN scramble_nonce_i[32] 
  END scramble_nonce_i[32]
  PIN scramble_nonce_i[31] 
  END scramble_nonce_i[31]
  PIN scramble_nonce_i[30] 
  END scramble_nonce_i[30]
  PIN scramble_nonce_i[29] 
  END scramble_nonce_i[29]
  PIN scramble_nonce_i[28] 
  END scramble_nonce_i[28]
  PIN scramble_nonce_i[27] 
  END scramble_nonce_i[27]
  PIN scramble_nonce_i[26] 
  END scramble_nonce_i[26]
  PIN scramble_nonce_i[25] 
  END scramble_nonce_i[25]
  PIN scramble_nonce_i[24] 
  END scramble_nonce_i[24]
  PIN scramble_nonce_i[23] 
  END scramble_nonce_i[23]
  PIN scramble_nonce_i[22] 
  END scramble_nonce_i[22]
  PIN scramble_nonce_i[21] 
  END scramble_nonce_i[21]
  PIN scramble_nonce_i[20] 
  END scramble_nonce_i[20]
  PIN scramble_nonce_i[19] 
  END scramble_nonce_i[19]
  PIN scramble_nonce_i[18] 
  END scramble_nonce_i[18]
  PIN scramble_nonce_i[17] 
  END scramble_nonce_i[17]
  PIN scramble_nonce_i[16] 
  END scramble_nonce_i[16]
  PIN scramble_nonce_i[15] 
  END scramble_nonce_i[15]
  PIN scramble_nonce_i[14] 
  END scramble_nonce_i[14]
  PIN scramble_nonce_i[13] 
  END scramble_nonce_i[13]
  PIN scramble_nonce_i[12] 
  END scramble_nonce_i[12]
  PIN scramble_nonce_i[11] 
  END scramble_nonce_i[11]
  PIN scramble_nonce_i[10] 
  END scramble_nonce_i[10]
  PIN scramble_nonce_i[9] 
  END scramble_nonce_i[9]
  PIN scramble_nonce_i[8] 
  END scramble_nonce_i[8]
  PIN scramble_nonce_i[7] 
  END scramble_nonce_i[7]
  PIN scramble_nonce_i[6] 
  END scramble_nonce_i[6]
  PIN scramble_nonce_i[5] 
  END scramble_nonce_i[5]
  PIN scramble_nonce_i[4] 
  END scramble_nonce_i[4]
  PIN scramble_nonce_i[3] 
  END scramble_nonce_i[3]
  PIN scramble_nonce_i[2] 
  END scramble_nonce_i[2]
  PIN scramble_nonce_i[1] 
  END scramble_nonce_i[1]
  PIN scramble_nonce_i[0] 
  END scramble_nonce_i[0]
  PIN debug_req_i 
    ANTENNAPARTIALMETALAREA 0.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.2477 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 112.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END debug_req_i
  PIN crash_dump_o[159] 
    ANTENNAPARTIALMETALAREA 5.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.054 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.97 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.02391 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 7.48943 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0538721 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 30.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 115.736 LAYER M3 ;
    ANTENNAGATEAREA 3.6684 LAYER M3 ; 
    ANTENNAMAXAREACAR 79.6025 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 307.987 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END crash_dump_o[159]
  PIN crash_dump_o[158] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 53.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 202.168 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.858 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.0228 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 137.004 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.41844 LAYER VL ;
  END crash_dump_o[158]
  PIN crash_dump_o[157] 
    ANTENNAPARTIALMETALAREA 4.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 28.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 105.672 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2972 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.7812 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 75.6895 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[157]
  PIN crash_dump_o[156] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.632 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.3692 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.2155 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.291 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[156]
  PIN crash_dump_o[155] 
    ANTENNAPARTIALMETALAREA 4.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 59.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 223.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.3692 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.6778 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 94.0604 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END crash_dump_o[155]
  PIN crash_dump_o[154] 
    ANTENNAPARTIALMETALAREA 1.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.29 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 48.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 180.264 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0016 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.0553 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.252 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.45098 LAYER VL ;
  END crash_dump_o[154]
  PIN crash_dump_o[153] 
    ANTENNAPARTIALMETALAREA 5.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.534 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 44.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 165.168 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.654 LAYER M3 ; 
    ANTENNAMAXAREACAR 47.1127 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 180.158 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END crash_dump_o[153]
  PIN crash_dump_o[152] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 52.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 196.544 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.654 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.601 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 143.617 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[152]
  PIN crash_dump_o[151] 
    ANTENNAPARTIALMETALAREA 0.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 45.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 168.72 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1364 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.1804 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 155.231 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END crash_dump_o[151]
  PIN crash_dump_o[150] 
    ANTENNAPARTIALMETALAREA 1.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.402 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 46.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 173.456 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.3692 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.5667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 96.2841 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.823045 LAYER VL ;
  END crash_dump_o[150]
  PIN crash_dump_o[149] 
    ANTENNAPARTIALMETALAREA 3.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.062 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 35.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 134.976 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.654 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.473 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 167.571 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END crash_dump_o[149]
  PIN crash_dump_o[148] 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 31.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 118.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9396 LAYER M3 ; 
    ANTENNAMAXAREACAR 157.604 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 589.94 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END crash_dump_o[148]
  PIN crash_dump_o[147] 
    ANTENNAPARTIALMETALAREA 6.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.162 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 36.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 138.232 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.3692 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.7289 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 94.2304 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.64609 LAYER VL ;
  END crash_dump_o[147]
  PIN crash_dump_o[146] 
    ANTENNAPARTIALMETALAREA 9.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.15 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.416 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.472 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.3195 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 141.83 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.41844 LAYER VL ;
  END crash_dump_o[146]
  PIN crash_dump_o[145] 
    ANTENNAPARTIALMETALAREA 5.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.462 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 101.232 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.86 LAYER M3 ; 
    ANTENNAMAXAREACAR 49.4329 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 194.227 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.44033 LAYER VL ;
  END crash_dump_o[145]
  PIN crash_dump_o[144] 
    ANTENNAPARTIALMETALAREA 9.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.706 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2972 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.0307 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 139.404 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.8018 LAYER VL ;
  END crash_dump_o[144]
  PIN crash_dump_o[143] 
    ANTENNAPARTIALMETALAREA 2.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.878 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 81.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.566 LAYER M3 ; 
    ANTENNAMAXAREACAR 80.4718 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 299.312 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[143]
  PIN crash_dump_o[142] 
    ANTENNAPARTIALMETALAREA 1.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.504 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2972 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.69997 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 29.3363 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[142]
  PIN crash_dump_o[141] 
    ANTENNAPARTIALMETALAREA 1.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.142 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 29.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 111.296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.5672 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.1796 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 63.6187 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[141]
  PIN crash_dump_o[140] 
    ANTENNAPARTIALMETALAREA 4.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.65 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.5672 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.6516 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 80.7715 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.23457 LAYER VL ;
  END crash_dump_o[140]
  PIN crash_dump_o[139] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2972 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.6912 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 82.95 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER VL ;
  END crash_dump_o[139]
  PIN crash_dump_o[138] 
    ANTENNAPARTIALMETALAREA 2.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.434 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 51 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 192.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.764 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.4452 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 145.253 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[138]
  PIN crash_dump_o[137] 
    ANTENNAPARTIALMETALAREA 3.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.062 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 31.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 118.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.9896 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.6331 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 100.67 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.408998 LAYER VL ;
  END crash_dump_o[137]
  PIN crash_dump_o[136] 
    ANTENNAPARTIALMETALAREA 11.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 43.216 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3996 LAYER M2 ; 
    ANTENNAMAXAREACAR 4.34246 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 16.5036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.116642 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 83.768 LAYER M3 ;
    ANTENNAGATEAREA 4.1364 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.0327 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 66.8046 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[136]
  PIN crash_dump_o[135] 
    ANTENNAPARTIALMETALAREA 8.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.822 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.52 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.658182 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2.23909 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER VL ;
  END crash_dump_o[135]
  PIN crash_dump_o[134] 
    ANTENNAPARTIALMETALAREA 9.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.594 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 83.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5752 LAYER M3 ; 
    ANTENNAMAXAREACAR 44.3468 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 171.376 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.64609 LAYER VL ;
  END crash_dump_o[134]
  PIN crash_dump_o[133] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 88.504 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6728 LAYER M3 ; 
    ANTENNAMAXAREACAR 55.5191 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 210.27 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.45098 LAYER VL ;
  END crash_dump_o[133]
  PIN crash_dump_o[132] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 29.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 114.552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8384 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.9657 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 115.291 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[132]
  PIN crash_dump_o[131] 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.52 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.906136 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.07239 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0227273 LAYER V2 ;
  END crash_dump_o[131]
  PIN crash_dump_o[130] 
    ANTENNAPARTIALMETALAREA 5.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.906 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.5456 LAYER M3 ; 
    ANTENNAMAXAREACAR 81.6912 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 304.712 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END crash_dump_o[130]
  PIN crash_dump_o[129] 
    ANTENNAPARTIALMETALAREA 3.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.766 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 28.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 109.224 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.024 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.1742 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 65.2312 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[129]
  PIN crash_dump_o[127] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 152.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 567.728 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.9896 LAYER M3 ; 
    ANTENNAMAXAREACAR 83.6619 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 313.859 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.77778 LAYER VL ;
  END crash_dump_o[127]
  PIN crash_dump_o[126] 
    ANTENNAPARTIALMETALAREA 3.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.618 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 36.9054 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 137.189 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.52 LAYER M3 ;
    ANTENNAGATEAREA 2.542 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.619 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 151.162 LAYER M3 ;
    ANTENNAMAXCUTCAR 5.55556 LAYER VL ;
  END crash_dump_o[126]
  PIN crash_dump_o[125] 
    ANTENNAPARTIALMETALAREA 3.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.726 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.32 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3664 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.7824 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 60.1514 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER VL ;
  END crash_dump_o[125]
  PIN crash_dump_o[124] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 42.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 158.064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2324 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.2896 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 88.6541 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[124]
  PIN crash_dump_o[123] 
    ANTENNAPARTIALMETALAREA 5.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 101.824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2324 LAYER M3 ; 
    ANTENNAMAXAREACAR 75.2588 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 285.095 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VL ;
  END crash_dump_o[123]
  PIN crash_dump_o[122] 
    ANTENNAPARTIALMETALAREA 3.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.098 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 45.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 173.16 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.4052 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.6655 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 121.03 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[122]
  PIN crash_dump_o[121] 
    ANTENNAPARTIALMETALAREA 1.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.402 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 37.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 140.896 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2324 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.3472 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 124.744 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.44174 LAYER VL ;
  END crash_dump_o[121]
  PIN crash_dump_o[120] 
    ANTENNAPARTIALMETALAREA 7.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.674 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 167.903 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 655.187 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAMAXCUTCAR 5.55556 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.272 LAYER M3 ;
    ANTENNAGATEAREA 4.2324 LAYER M3 ; 
    ANTENNAMAXAREACAR 171.608 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 669.664 LAYER M3 ;
    ANTENNAMAXCUTCAR 5.55556 LAYER VL ;
  END crash_dump_o[120]
  PIN crash_dump_o[119] 
    ANTENNAPARTIALMETALAREA 1.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 80.216 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2324 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.4907 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 75.689 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.77778 LAYER VL ;
  END crash_dump_o[119]
  PIN crash_dump_o[118] 
    ANTENNAPARTIALMETALAREA 4.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 74.592 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1104 LAYER M3 ; 
    ANTENNAMAXAREACAR 64.0156 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 248.286 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VL ;
  END crash_dump_o[118]
  PIN crash_dump_o[117] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.47 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 35.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 134.68 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2324 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.7977 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.571 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.56341 LAYER VL ;
  END crash_dump_o[117]
  PIN crash_dump_o[116] 
    ANTENNAPARTIALMETALAREA 5.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.682 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 31.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 121.656 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2324 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.2824 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 55.0773 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[116]
  PIN crash_dump_o[115] 
    ANTENNAPARTIALMETALAREA 5.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.87 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.544 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1104 LAYER M3 ; 
    ANTENNAMAXAREACAR 53.5806 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 202.157 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[115]
  PIN crash_dump_o[114] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.304 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.962 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.39014 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 26.2492 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END crash_dump_o[114]
  PIN crash_dump_o[113] 
    ANTENNAPARTIALMETALAREA 9.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 36.778 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.848 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.91847 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 14.6041 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0561798 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 56.24 LAYER M3 ;
    ANTENNAGATEAREA 3.1936 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.5986 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 86.0477 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[113]
  PIN crash_dump_o[112] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.24 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.962 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.0709 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 69.5181 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END crash_dump_o[112]
  PIN crash_dump_o[111] 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.622 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.608 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4548 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.1848 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.317 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VL ;
  END crash_dump_o[111]
  PIN crash_dump_o[110] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.32 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2324 LAYER M3 ; 
    ANTENNAMAXAREACAR 52.8865 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 197.528 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.77778 LAYER VL ;
  END crash_dump_o[110]
  PIN crash_dump_o[109] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.512 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1104 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.1193 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 188.653 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[109]
  PIN crash_dump_o[108] 
    ANTENNAPARTIALMETALAREA 6.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.05 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.568 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2324 LAYER M3 ; 
    ANTENNAMAXAREACAR 146.906 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 546.911 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.77778 LAYER VL ;
  END crash_dump_o[108]
  PIN crash_dump_o[107] 
    ANTENNAPARTIALMETALAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.838 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.014 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.31102 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 8.72115 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0595829 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.92 LAYER M3 ;
    ANTENNAGATEAREA 2.962 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.09876 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 25.0212 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[107]
  PIN crash_dump_o[106] 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.698 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.144 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1748 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.00406 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 34.403 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.746269 LAYER VL ;
  END crash_dump_o[106]
  PIN crash_dump_o[105] 
    ANTENNAPARTIALMETALAREA 3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.396 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.97 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.24949 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 4.57428 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.040404 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 52.392 LAYER M3 ;
    ANTENNAGATEAREA 4.2324 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.5177 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 124.754 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VL ;
  END crash_dump_o[105]
  PIN crash_dump_o[104] 
    ANTENNAPARTIALMETALAREA 4.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.946 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 78.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 295.408 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2324 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.7477 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 101.269 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.77778 LAYER VL ;
  END crash_dump_o[104]
  PIN crash_dump_o[103] 
    ANTENNAPARTIALMETALAREA 7.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.64 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.848 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.16032 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 11.9374 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0842697 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.144 LAYER M3 ;
    ANTENNAGATEAREA 3.3328 LAYER M3 ; 
    ANTENNAMAXAREACAR 68.3796 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 257.218 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VL ;
  END crash_dump_o[103]
  PIN crash_dump_o[102] 
    ANTENNAPARTIALMETALAREA 11.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 41.514 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 41.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 154.808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1104 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.2317 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 120.762 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[102]
  PIN crash_dump_o[101] 
    ANTENNAPARTIALMETALAREA 2.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.99 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 87.024 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5152 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.4987 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 151.611 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END crash_dump_o[101]
  PIN crash_dump_o[100] 
    ANTENNAPARTIALMETALAREA 6.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.754 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.048 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4644 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.3994 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 69.7838 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.83062 LAYER VL ;
  END crash_dump_o[100]
  PIN crash_dump_o[99] 
    ANTENNAPARTIALMETALAREA 8.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.414 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4068 LAYER M3 ; 
    ANTENNAMAXAREACAR 114.707 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 425.289 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.394605 LAYER VL ;
  END crash_dump_o[99]
  PIN crash_dump_o[98] 
    ANTENNAPARTIALMETALAREA 1.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 43.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 166.352 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4644 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.8881 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 90.3966 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[98]
  PIN crash_dump_o[97] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 34.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 126.392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8744 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.3425 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 70.3275 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[97]
  PIN crash_dump_o[95] 
    ANTENNAPARTIALMETALAREA 9.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.558 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.008 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2152 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.40572 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 17.5059 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[95]
  PIN crash_dump_o[94] 
    ANTENNAPARTIALMETALAREA 7.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.378 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1128 LAYER M2 ; 
    ANTENNAMAXAREACAR 70.4894 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 264.181 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.408 LAYER M3 ;
    ANTENNAGATEAREA 3.8272 LAYER M3 ; 
    ANTENNAMAXAREACAR 73.0291 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 273.694 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER VL ;
  END crash_dump_o[94]
  PIN crash_dump_o[93] 
    ANTENNAPARTIALMETALAREA 3.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.766 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.112 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9088 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.63122 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 18.2325 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.411523 LAYER VL ;
  END crash_dump_o[93]
  PIN crash_dump_o[92] 
    ANTENNAPARTIALMETALAREA 2.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8272 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.5537 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 59.5889 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER VL ;
  END crash_dump_o[92]
  PIN crash_dump_o[91] 
    ANTENNAPARTIALMETALAREA 3.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.726 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 59.2 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8272 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.3043 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 140.182 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER VL ;
  END crash_dump_o[91]
  PIN crash_dump_o[90] 
    ANTENNAPARTIALMETALAREA 3.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.098 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.616 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.024 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.3562 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 40.281 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.41844 LAYER VL ;
  END crash_dump_o[90]
  PIN crash_dump_o[89] 
    ANTENNAPARTIALMETALAREA 3.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.062 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.32 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9088 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.0838 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 100.714 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02881 LAYER VL ;
  END crash_dump_o[89]
  PIN crash_dump_o[88] 
    ANTENNAPARTIALMETALAREA 15.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.682 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 LAYER M2 ; 
    ANTENNAMAXAREACAR 82.3807 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 304.626 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.617284 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.24 LAYER M3 ;
    ANTENNAGATEAREA 3.9088 LAYER M3 ; 
    ANTENNAMAXAREACAR 83.6394 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 309.548 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.617284 LAYER VL ;
  END crash_dump_o[88]
  PIN crash_dump_o[87] 
    ANTENNAPARTIALMETALAREA 15.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.238 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.672 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1056 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.5684 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 44.7604 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.823045 LAYER VL ;
  END crash_dump_o[87]
  PIN crash_dump_o[86] 
    ANTENNAPARTIALMETALAREA 3.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.506 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.72 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8272 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.40423 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 21.6976 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER VL ;
  END crash_dump_o[86]
  PIN crash_dump_o[85] 
    ANTENNAPARTIALMETALAREA 10.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 38.702 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.048 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8272 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.1993 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 91.3167 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.77305 LAYER VL ;
  END crash_dump_o[85]
  PIN crash_dump_o[84] 
    ANTENNAPARTIALMETALAREA 14.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 52.466 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8272 LAYER M3 ; 
    ANTENNAMAXAREACAR 69.8544 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 270.36 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER VL ;
  END crash_dump_o[84]
  PIN crash_dump_o[83] 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.214 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.92 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8272 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.2343 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 104.684 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.875443 LAYER VL ;
  END crash_dump_o[83]
  PIN crash_dump_o[82] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7456 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.8809 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 46.7718 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END crash_dump_o[82]
  PIN crash_dump_o[81] 
    ANTENNAPARTIALMETALAREA 10.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 39.59 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.464 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8272 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.7622 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 48.8833 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER VL ;
  END crash_dump_o[81]
  PIN crash_dump_o[80] 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.698 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.52 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8272 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.0813 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 46.5575 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.41844 LAYER VL ;
  END crash_dump_o[80]
  PIN crash_dump_o[79] 
    ANTENNAPARTIALMETALAREA 6.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.902 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3912 LAYER M2 ; 
    ANTENNAMAXAREACAR 18.6104 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 69.8425 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.613497 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.144 LAYER M3 ;
    ANTENNAGATEAREA 4.084 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.8723 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.5721 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[79]
  PIN crash_dump_o[78] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.568 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.7136 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 131.503 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[78]
  PIN crash_dump_o[77] 
    ANTENNAPARTIALMETALAREA 3.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.766 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.936 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.3726 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 141.816 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[77]
  PIN crash_dump_o[76] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.464 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.9188 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 118.958 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[76]
  PIN crash_dump_o[75] 
    ANTENNAPARTIALMETALAREA 4.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.13 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.704 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.8892 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 52.8427 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[75]
  PIN crash_dump_o[74] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.784 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.084 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.6377 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 43.0724 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[74]
  PIN crash_dump_o[73] 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.084 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.0257 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.6393 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[73]
  PIN crash_dump_o[72] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.016 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.084 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.81021 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 37.3284 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[72]
  PIN crash_dump_o[71] 
    ANTENNAPARTIALMETALAREA 1.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.958 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 78.144 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.8056 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 90.0021 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[71]
  PIN crash_dump_o[70] 
    ANTENNAPARTIALMETALAREA 1.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.474 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 74.888 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.6747 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 141.92 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VL ;
  END crash_dump_o[70]
  PIN crash_dump_o[69] 
    ANTENNAPARTIALMETALAREA 10.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 39.294 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 74.296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.784 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.948 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 43.6802 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.29885 LAYER VL ;
  END crash_dump_o[69]
  PIN crash_dump_o[68] 
    ANTENNAPARTIALMETALAREA 2.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.73 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 96.792 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8248 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.8134 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 134.855 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.51515 LAYER VL ;
  END crash_dump_o[68]
  PIN crash_dump_o[67] 
    ANTENNAPARTIALMETALAREA 4.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.428 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 33.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 124.912 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8248 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.8909 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 80.5404 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.909091 LAYER VL ;
  END crash_dump_o[67]
  PIN crash_dump_o[66] 
    ANTENNAPARTIALMETALAREA 15.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 57.498 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 89.392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.288 LAYER M3 ; 
    ANTENNAMAXAREACAR 60.1481 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 232.019 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.87356 LAYER VL ;
  END crash_dump_o[66]
  PIN crash_dump_o[65] 
    ANTENNAPARTIALMETALAREA 27.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 104.414 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 104.192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9976 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.48116 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 36.5 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.909091 LAYER VL ;
  END crash_dump_o[65]
  PIN crash_dump_o[64] 
    ANTENNAPARTIALMETALAREA 2.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.138 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 81.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 305.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.024 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.5775 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 113.217 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END crash_dump_o[64]
  PIN crash_dump_o[63] 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.214 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 46.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 176.12 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3612 LAYER M3 ; 
    ANTENNAMAXAREACAR 58.3811 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 226.915 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.5977 LAYER VL ;
  END crash_dump_o[63]
  PIN crash_dump_o[62] 
    ANTENNAPARTIALMETALAREA 9.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.002 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 34.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 130.832 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.27 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.5021 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 92.3891 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.29885 LAYER VL ;
  END crash_dump_o[62]
  PIN crash_dump_o[61] 
    ANTENNAPARTIALMETALAREA 6.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.974 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 55.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 208.088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4428 LAYER M3 ; 
    ANTENNAMAXAREACAR 70.034 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 268.414 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[61]
  PIN crash_dump_o[60] 
    ANTENNAPARTIALMETALAREA 3.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.21 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 42.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 163.096 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4428 LAYER M3 ; 
    ANTENNAMAXAREACAR 68.016 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 272.35 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.5977 LAYER VL ;
  END crash_dump_o[60]
  PIN crash_dump_o[59] 
    ANTENNAPARTIALMETALAREA 8.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.19 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 122.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4 LAYER M3 ; 
    ANTENNAMAXAREACAR 132.152 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 506.185 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[59]
  PIN crash_dump_o[58] 
    ANTENNAPARTIALMETALAREA 2.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.434 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.148 LAYER M3 ; 
    ANTENNAMAXAREACAR 147.875 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 551.623 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.29885 LAYER VL ;
  END crash_dump_o[58]
  PIN crash_dump_o[57] 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 28.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 110.112 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.148 LAYER M3 ; 
    ANTENNAMAXAREACAR 52.0909 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 210.162 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.5977 LAYER VL ;
  END crash_dump_o[57]
  PIN crash_dump_o[56] 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.16 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.148 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.818 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 182.539 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.5977 LAYER VL ;
  END crash_dump_o[56]
  PIN crash_dump_o[55] 
    ANTENNAPARTIALMETALAREA 3.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.654 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 34.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 131.128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.148 LAYER M3 ; 
    ANTENNAMAXAREACAR 62.2038 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 251.275 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[55]
  PIN crash_dump_o[54] 
    ANTENNAPARTIALMETALAREA 4.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.538 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 75.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 282.976 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4428 LAYER M3 ; 
    ANTENNAMAXAREACAR 65.119 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 254.113 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.29885 LAYER VL ;
  END crash_dump_o[54]
  PIN crash_dump_o[53] 
    ANTENNAPARTIALMETALAREA 11.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 40.774 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 38.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 145.928 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.27 LAYER M3 ; 
    ANTENNAMAXAREACAR 44.828 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 173.557 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.02299 LAYER VL ;
  END crash_dump_o[53]
  PIN crash_dump_o[52] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 82.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.27 LAYER M3 ; 
    ANTENNAMAXAREACAR 63.8813 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 241.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.87356 LAYER VL ;
  END crash_dump_o[52]
  PIN crash_dump_o[51] 
    ANTENNAPARTIALMETALAREA 16.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.198 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 63.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 237.096 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.27 LAYER M3 ; 
    ANTENNAMAXAREACAR 87.2887 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 337.713 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.5977 LAYER VL ;
  END crash_dump_o[51]
  PIN crash_dump_o[50] 
    ANTENNAPARTIALMETALAREA 2.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.026 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 88.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 330.336 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2124 LAYER M3 ; 
    ANTENNAMAXAREACAR 51.3752 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 194.521 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.44828 LAYER VL ;
  END crash_dump_o[50]
  PIN crash_dump_o[49] 
    ANTENNAPARTIALMETALAREA 10.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 40.182 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 47.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 180.264 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4428 LAYER M3 ; 
    ANTENNAMAXAREACAR 43.7868 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 171.686 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[49]
  PIN crash_dump_o[48] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 50 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 188.256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4428 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.7745 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.187 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.29885 LAYER VL ;
  END crash_dump_o[48]
  PIN crash_dump_o[47] 
    ANTENNAPARTIALMETALAREA 10.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 39.886 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 123.432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.27 LAYER M3 ; 
    ANTENNAMAXAREACAR 129.839 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 497.525 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[47]
  PIN crash_dump_o[46] 
    ANTENNAPARTIALMETALAREA 5.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.386 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 52.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 197.432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.27 LAYER M3 ; 
    ANTENNAMAXAREACAR 61.6919 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 241.676 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.5977 LAYER VL ;
  END crash_dump_o[46]
  PIN crash_dump_o[45] 
    ANTENNAPARTIALMETALAREA 1.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 61.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 234.432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.27 LAYER M3 ; 
    ANTENNAMAXAREACAR 87.9292 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 339.933 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[45]
  PIN crash_dump_o[44] 
    ANTENNAPARTIALMETALAREA 4.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.834 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 51.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 193.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.27 LAYER M3 ; 
    ANTENNAMAXAREACAR 102.938 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 395.644 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[44]
  PIN crash_dump_o[43] 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.25 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 58.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 222.592 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.27 LAYER M3 ; 
    ANTENNAMAXAREACAR 55.0485 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 206.383 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.29885 LAYER VL ;
  END crash_dump_o[43]
  PIN crash_dump_o[42] 
    ANTENNAPARTIALMETALAREA 3.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.506 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 69.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 264.92 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3324 LAYER M3 ; 
    ANTENNAMAXAREACAR 44.0954 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 169.276 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[42]
  PIN crash_dump_o[41] 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.214 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 51.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 194.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.27 LAYER M3 ; 
    ANTENNAMAXAREACAR 55.4859 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 211.194 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.87356 LAYER VL ;
  END crash_dump_o[41]
  PIN crash_dump_o[40] 
    ANTENNAPARTIALMETALAREA 5.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.314 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 29.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 114.256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3324 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.9276 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 99.4712 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.42424 LAYER VL ;
  END crash_dump_o[40]
  PIN crash_dump_o[39] 
    ANTENNAPARTIALMETALAREA 0.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.478 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 45.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 168.424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.834 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.4485 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 151.192 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[39]
  PIN crash_dump_o[38] 
    ANTENNAPARTIALMETALAREA 23.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 87.098 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 50.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 189.144 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4428 LAYER M3 ; 
    ANTENNAMAXAREACAR 119.959 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 458.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[38]
  PIN crash_dump_o[37] 
    ANTENNAPARTIALMETALAREA 5.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.126 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 39.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 150.96 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7956 LAYER M3 ; 
    ANTENNAMAXAREACAR 53.0922 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 204.163 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[37]
  PIN crash_dump_o[36] 
    ANTENNAPARTIALMETALAREA 6.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.754 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 43.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 167.536 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.27 LAYER M3 ; 
    ANTENNAMAXAREACAR 66.9254 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 262.407 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[36]
  PIN crash_dump_o[35] 
    ANTENNAPARTIALMETALAREA 5.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 72.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 273.208 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3732 LAYER M3 ; 
    ANTENNAMAXAREACAR 49.713 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 191.327 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[35]
  PIN crash_dump_o[34] 
    ANTENNAPARTIALMETALAREA 3.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.098 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 66.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 248.048 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.546 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.3665 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 88.848 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.73408 LAYER VL ;
  END crash_dump_o[34]
  PIN crash_dump_o[33] 
    ANTENNAPARTIALMETALAREA 1.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.07 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 93.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 351.944 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3132 LAYER M3 ; 
    ANTENNAMAXAREACAR 69.5272 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 262.808 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.77778 LAYER VL ;
  END crash_dump_o[33]
  PIN crash_dump_o[32] 
    ANTENNAPARTIALMETALAREA 3.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.21 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 50.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 192.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2004 LAYER M3 ; 
    ANTENNAMAXAREACAR 107.929 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 417.21 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.47222 LAYER VL ;
  END crash_dump_o[32]
  PIN crash_dump_o[31] 
    ANTENNAPARTIALMETALAREA 24.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 92.574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 59.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 221.408 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.9374 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 82.0025 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[31]
  PIN crash_dump_o[30] 
    ANTENNAPARTIALMETALAREA 48.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 181.226 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 100.344 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.8308 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 59.0194 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[30]
  PIN crash_dump_o[29] 
    ANTENNAPARTIALMETALAREA 3.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.654 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 100.64 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1936 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.3941 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 51.116 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[29]
  PIN crash_dump_o[28] 
    ANTENNAPARTIALMETALAREA 41.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 155.474 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 37.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 137.936 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1936 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.613 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 81.8453 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[28]
  PIN crash_dump_o[27] 
    ANTENNAPARTIALMETALAREA 39.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 145.262 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.6 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1936 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.21268 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 32.0405 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[27]
  PIN crash_dump_o[26] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 34.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 132.016 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0208 LAYER M3 ; 
    ANTENNAMAXAREACAR 63.452 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 245.575 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[26]
  PIN crash_dump_o[25] 
    ANTENNAPARTIALMETALAREA 3.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.062 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 70.448 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0208 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.2004 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 46.4853 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[25]
  PIN crash_dump_o[24] 
    ANTENNAPARTIALMETALAREA 1.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.474 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 50.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 190.328 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0208 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.8727 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 89.9757 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[24]
  PIN crash_dump_o[23] 
    ANTENNAPARTIALMETALAREA 6.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.79 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 52.984 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0208 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.7965 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 44.5096 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[23]
  PIN crash_dump_o[22] 
    ANTENNAPARTIALMETALAREA 6.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.866 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1936 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.1401 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 38.4926 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[22]
  PIN crash_dump_o[21] 
    ANTENNAPARTIALMETALAREA 20.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 77.182 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 45.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 170.2 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.058 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 67.8338 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[21]
  PIN crash_dump_o[20] 
    ANTENNAPARTIALMETALAREA 10.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 37.962 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 36.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 137.344 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.5114 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 62.0044 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[20]
  PIN crash_dump_o[19] 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.102 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 108.04 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0208 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.4433 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 141.532 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[19]
  PIN crash_dump_o[18] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 52.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 196.248 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0208 LAYER M3 ; 
    ANTENNAMAXAREACAR 48.7625 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 186.607 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[18]
  PIN crash_dump_o[17] 
    ANTENNAPARTIALMETALAREA 8.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.822 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 46.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 175.232 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3156 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.5684 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 139.928 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[17]
  PIN crash_dump_o[16] 
    ANTENNAPARTIALMETALAREA 5.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.57 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 79.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3156 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.6662 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 119.364 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[16]
  PIN crash_dump_o[15] 
    ANTENNAPARTIALMETALAREA 5.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.534 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 43.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 161.024 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.939 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 170.604 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[15]
  PIN crash_dump_o[14] 
    ANTENNAPARTIALMETALAREA 8.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.226 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 51.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 192.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.3919 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 172.303 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[14]
  PIN crash_dump_o[13] 
    ANTENNAPARTIALMETALAREA 44.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 163.91 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 29.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 114.552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.9588 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 76.5625 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[13]
  PIN crash_dump_o[12] 
    ANTENNAPARTIALMETALAREA 9.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 36.186 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 56.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 214.008 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0372 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.2501 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.0337 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.19048 LAYER VL ;
  END crash_dump_o[12]
  PIN crash_dump_o[11] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.806 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 89.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 338.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.3731 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 125.963 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[11]
  PIN crash_dump_o[10] 
    ANTENNAPARTIALMETALAREA 17.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 66.378 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 43.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 164.872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.8858 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 67.7798 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[10]
  PIN crash_dump_o[9] 
    ANTENNAPARTIALMETALAREA 5.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.462 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 68.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 260.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.4191 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 96.1847 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[9]
  PIN crash_dump_o[8] 
    ANTENNAPARTIALMETALAREA 4.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.466 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 66.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 252.488 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 81.7376 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 312.864 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[8]
  PIN crash_dump_o[7] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.806 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 52.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 196.544 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6684 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.8588 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 78.4648 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.171821 LAYER VL ;
  END crash_dump_o[7]
  PIN crash_dump_o[6] 
    ANTENNAPARTIALMETALAREA 9.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 36.778 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 47.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 177.896 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3156 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.2439 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 73.0489 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER VL ;
  END crash_dump_o[6]
  PIN crash_dump_o[5] 
    ANTENNAPARTIALMETALAREA 8.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.19 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 42.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 158.656 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6684 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.0274 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 60.0839 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.171821 LAYER VL ;
  END crash_dump_o[5]
  PIN crash_dump_o[4] 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.698 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 42.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 161.32 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.8858 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 78.2999 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[4]
  PIN crash_dump_o[3] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.806 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 86.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 323.528 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.885 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 141.903 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[3]
  PIN crash_dump_o[2] 
    ANTENNAPARTIALMETALAREA 65.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 240.722 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 47.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 176.12 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3156 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.6696 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 66.2285 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER VL ;
  END crash_dump_o[2]
  PIN crash_dump_o[1] 
    ANTENNAPARTIALMETALAREA 51.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 191.438 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 82.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 309.024 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.501 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 128.723 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[1]
  PIN crash_dump_o[0] 
    ANTENNAPARTIALMETALAREA 51.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 190.698 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 63.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 237.688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1428 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.9662 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 86.267 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[0]
  PIN double_fault_seen_o 
    ANTENNAPARTIALMETALAREA 8.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 101.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 377.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.126 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.6931 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 125.281 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.282002 LAYER VL ;
  END double_fault_seen_o
  PIN fetch_enable_i[3] 
  END fetch_enable_i[3]
  PIN fetch_enable_i[2] 
  END fetch_enable_i[2]
  PIN fetch_enable_i[1] 
  END fetch_enable_i[1]
  PIN fetch_enable_i[0] 
  END fetch_enable_i[0]
  PIN core_sleep_o 
    ANTENNAPARTIALMETALAREA 0.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 35.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 132.608 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.98 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.9121 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 60.0599 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.21212 LAYER VL ;
  END core_sleep_o
  PIN scan_rst_ni 
  END scan_rst_ni
END ibex_top

END LIBRARY
