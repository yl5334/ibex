/courses/ee6321/share/ibm13rflpvt/lef/ibm13rflpvt_macros.lef