

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO ibex_top 
  PIN clk_i 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.208 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5976 LAYER M3 ; 
    ANTENNAMAXAREACAR 67.0509 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 249.814 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END clk_i
  PIN rst_ni 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.9369 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.329 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END rst_ni
  PIN test_en_i 
    ANTENNAPARTIALMETALAREA 1.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.6171 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END test_en_i
  PIN ram_cfg_i[9] 
  END ram_cfg_i[9]
  PIN ram_cfg_i[8] 
  END ram_cfg_i[8]
  PIN ram_cfg_i[7] 
  END ram_cfg_i[7]
  PIN ram_cfg_i[6] 
  END ram_cfg_i[6]
  PIN ram_cfg_i[5] 
  END ram_cfg_i[5]
  PIN ram_cfg_i[4] 
  END ram_cfg_i[4]
  PIN ram_cfg_i[3] 
  END ram_cfg_i[3]
  PIN ram_cfg_i[2] 
  END ram_cfg_i[2]
  PIN ram_cfg_i[1] 
  END ram_cfg_i[1]
  PIN ram_cfg_i[0] 
  END ram_cfg_i[0]
  PIN hart_id_i[31] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.7162 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 89.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[31]
  PIN hart_id_i[30] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.4414 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 119.995 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[30]
  PIN hart_id_i[29] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.6171 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[29]
  PIN hart_id_i[28] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.4189 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 99.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[28]
  PIN hart_id_i[27] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.4189 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 99.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[27]
  PIN hart_id_i[26] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.5856 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 99.9955 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[26]
  PIN hart_id_i[25] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.6171 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[25]
  PIN hart_id_i[24] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.1351 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 96.6622 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[24]
  PIN hart_id_i[23] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.7387 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.995 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[23]
  PIN hart_id_i[22] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.6171 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[22]
  PIN hart_id_i[21] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.1667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 89.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[21]
  PIN hart_id_i[20] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
  END hart_id_i[20]
  PIN hart_id_i[19] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.3198 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[19]
  PIN hart_id_i[18] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.3333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 89.9955 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[18]
  PIN hart_id_i[17] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
  END hart_id_i[17]
  PIN hart_id_i[16] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
  END hart_id_i[16]
  PIN hart_id_i[15] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.2342 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.3288 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[15]
  PIN hart_id_i[14] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
  END hart_id_i[14]
  PIN hart_id_i[13] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
  END hart_id_i[13]
  PIN hart_id_i[12] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3 ;
  END hart_id_i[12]
  PIN hart_id_i[11] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
  END hart_id_i[11]
  PIN hart_id_i[10] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.3198 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[10]
  PIN hart_id_i[9] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
  END hart_id_i[9]
  PIN hart_id_i[8] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
  END hart_id_i[8]
  PIN hart_id_i[7] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M3 ;
  END hart_id_i[7]
  PIN hart_id_i[6] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3 ;
  END hart_id_i[6]
  PIN hart_id_i[5] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
  END hart_id_i[5]
  PIN hart_id_i[4] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
  END hart_id_i[4]
  PIN hart_id_i[3] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
  END hart_id_i[3]
  PIN hart_id_i[2] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
  END hart_id_i[2]
  PIN hart_id_i[1] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.7838 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.3288 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[1]
  PIN hart_id_i[0] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.7162 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 89.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END hart_id_i[0]
  PIN boot_addr_i[31] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.92 LAYER M3 ;
  END boot_addr_i[31]
  PIN boot_addr_i[30] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
  END boot_addr_i[30]
  PIN boot_addr_i[29] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.1306 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 143.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END boot_addr_i[29]
  PIN boot_addr_i[28] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.8378 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 106.662 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END boot_addr_i[28]
  PIN boot_addr_i[27] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
  END boot_addr_i[27]
  PIN boot_addr_i[26] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.504 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.6892 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 173.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END boot_addr_i[26]
  PIN boot_addr_i[25] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.2883 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.995 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END boot_addr_i[25]
  PIN boot_addr_i[24] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.1306 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 143.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END boot_addr_i[24]
  PIN boot_addr_i[23] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.3874 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 106.662 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END boot_addr_i[23]
  PIN boot_addr_i[22] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.9459 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 136.662 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END boot_addr_i[22]
  PIN boot_addr_i[21] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER M3 ;
  END boot_addr_i[21]
  PIN boot_addr_i[20] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
  END boot_addr_i[20]
  PIN boot_addr_i[19] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.3198 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END boot_addr_i[19]
  PIN boot_addr_i[18] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.3198 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END boot_addr_i[18]
  PIN boot_addr_i[17] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
  END boot_addr_i[17]
  PIN boot_addr_i[16] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
  END boot_addr_i[16]
  PIN boot_addr_i[15] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
  END boot_addr_i[15]
  PIN boot_addr_i[14] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.4324 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 86.6622 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END boot_addr_i[14]
  PIN boot_addr_i[13] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.4324 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 86.6622 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END boot_addr_i[13]
  PIN boot_addr_i[12] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
  END boot_addr_i[12]
  PIN boot_addr_i[11] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
  END boot_addr_i[11]
  PIN boot_addr_i[10] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
  END boot_addr_i[10]
  PIN boot_addr_i[9] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
  END boot_addr_i[9]
  PIN boot_addr_i[8] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
  END boot_addr_i[8]
  PIN boot_addr_i[7] 
  END boot_addr_i[7]
  PIN boot_addr_i[6] 
  END boot_addr_i[6]
  PIN boot_addr_i[5] 
  END boot_addr_i[5]
  PIN boot_addr_i[4] 
  END boot_addr_i[4]
  PIN boot_addr_i[3] 
  END boot_addr_i[3]
  PIN boot_addr_i[2] 
  END boot_addr_i[2]
  PIN boot_addr_i[1] 
  END boot_addr_i[1]
  PIN boot_addr_i[0] 
  END boot_addr_i[0]
  PIN instr_req_o 
    ANTENNAPARTIALMETALAREA 8.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.56 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3 LAYER M3 ; 
    ANTENNAMAXAREACAR 158.209 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 586.476 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END instr_req_o
  PIN instr_gnt_i 
    ANTENNAPARTIALMETALAREA 2.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.508 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0696 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.9195 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 177.069 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.14943 LAYER VL ;
  END instr_gnt_i
  PIN instr_rvalid_i 
    ANTENNAPARTIALMETALAREA 2.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.2883 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 109.995 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_rvalid_i
  PIN instr_addr_o[31] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.14141 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.17125 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[31]
  PIN instr_addr_o[30] 
    ANTENNAPARTIALMETALAREA 3.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.54672 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.81891 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[30]
  PIN instr_addr_o[29] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.17266 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.28688 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[29]
  PIN instr_addr_o[28] 
    ANTENNAPARTIALMETALAREA 2.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.916 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.30453 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.92281 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[28]
  PIN instr_addr_o[27] 
    ANTENNAPARTIALMETALAREA 5.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.536 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.09359 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 11.34 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[27]
  PIN instr_addr_o[26] 
    ANTENNAPARTIALMETALAREA 6.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.124 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.77422 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 10.3572 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[26]
  PIN instr_addr_o[25] 
    ANTENNAPARTIALMETALAREA 5.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.904 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.57891 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.49 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[25]
  PIN instr_addr_o[24] 
    ANTENNAPARTIALMETALAREA 5.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.164 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.46172 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.20094 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[24]
  PIN instr_addr_o[23] 
    ANTENNAPARTIALMETALAREA 6.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.792 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.67266 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.83688 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[23]
  PIN instr_addr_o[22] 
    ANTENNAPARTIALMETALAREA 6.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.644 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.61797 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.77906 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[22]
  PIN instr_addr_o[21] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.066 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.70657 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.87054 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0750469 LAYER VL ;
  END instr_addr_o[21]
  PIN instr_addr_o[20] 
    ANTENNAPARTIALMETALAREA 2.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.916 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.30453 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.92281 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[20]
  PIN instr_addr_o[19] 
    ANTENNAPARTIALMETALAREA 2.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.656 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.39141 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.09625 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[19]
  PIN instr_addr_o[18] 
    ANTENNAPARTIALMETALAREA 2.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.14 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.08672 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.11344 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[18]
  PIN instr_addr_o[17] 
    ANTENNAPARTIALMETALAREA 5.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.312 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.51641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.25875 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[17]
  PIN instr_addr_o[16] 
    ANTENNAPARTIALMETALAREA 6.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.94 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.64922 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.89469 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[16]
  PIN instr_addr_o[15] 
    ANTENNAPARTIALMETALAREA 5.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.72 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.48422 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.14312 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[15]
  PIN instr_addr_o[14] 
    ANTENNAPARTIALMETALAREA 5.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.682 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.50078 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.40328 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[14]
  PIN instr_addr_o[13] 
    ANTENNAPARTIALMETALAREA 4.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.984 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.95391 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.1775 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[13]
  PIN instr_addr_o[12] 
    ANTENNAPARTIALMETALAREA 2.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.14 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.11703 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.22906 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[12]
  PIN instr_addr_o[11] 
    ANTENNAPARTIALMETALAREA 5.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.24 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.29766 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.44937 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[11]
  PIN instr_addr_o[10] 
    ANTENNAPARTIALMETALAREA 3.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.06 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.10141 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 15.2134 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[10]
  PIN instr_addr_o[9] 
    ANTENNAPARTIALMETALAREA 5.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.56234 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 16.7744 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[9]
  PIN instr_addr_o[8] 
    ANTENNAPARTIALMETALAREA 4.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.132 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.96078 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.35094 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[8]
  PIN instr_addr_o[7] 
    ANTENNAPARTIALMETALAREA 5.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.944 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.26641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.33375 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.03125 LAYER VL ;
  END instr_addr_o[7]
  PIN instr_addr_o[6] 
    ANTENNAPARTIALMETALAREA 4.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.316 LAYER M3 ;
  END instr_addr_o[6]
  PIN instr_addr_o[5] 
    ANTENNAPARTIALMETALAREA 3.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.024 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.17109 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.25816 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0197824 LAYER VL ;
  END instr_addr_o[5]
  PIN instr_addr_o[4] 
    ANTENNAPARTIALMETALAREA 3.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.356 LAYER M3 ;
  END instr_addr_o[4]
  PIN instr_addr_o[3] 
    ANTENNAPARTIALMETALAREA 4.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.168 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.43301 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.21978 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0197824 LAYER VL ;
  END instr_addr_o[3]
  PIN instr_addr_o[2] 
    ANTENNAPARTIALMETALAREA 5.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.388 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.044 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.55665 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.76874 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0197824 LAYER VL ;
  END instr_addr_o[2]
  PIN instr_rdata_i[31] 
    ANTENNAPARTIALMETALAREA 1.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
  END instr_rdata_i[31]
  PIN instr_rdata_i[30] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M3 ;
  END instr_rdata_i[30]
  PIN instr_rdata_i[29] 
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.512 LAYER M3 ;
  END instr_rdata_i[29]
  PIN instr_rdata_i[28] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M3 ;
  END instr_rdata_i[28]
  PIN instr_rdata_i[27] 
    ANTENNAPARTIALMETALAREA 0.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
  END instr_rdata_i[27]
  PIN instr_rdata_i[26] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M3 ;
  END instr_rdata_i[26]
  PIN instr_rdata_i[25] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.3333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 89.9955 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_rdata_i[25]
  PIN instr_rdata_i[24] 
    ANTENNAPARTIALMETALAREA 1.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.364 LAYER M3 ;
  END instr_rdata_i[24]
  PIN instr_rdata_i[23] 
    ANTENNAPARTIALMETALAREA 2.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.1892 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 113.329 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_rdata_i[23]
  PIN instr_rdata_i[22] 
    ANTENNAPARTIALMETALAREA 1.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.364 LAYER M3 ;
  END instr_rdata_i[22]
  PIN instr_rdata_i[21] 
    ANTENNAPARTIALMETALAREA 2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.518 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 96.3559 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_rdata_i[21]
  PIN instr_rdata_i[20] 
    ANTENNAPARTIALMETALAREA 1.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.66 LAYER M3 ;
  END instr_rdata_i[20]
  PIN instr_rdata_i[19] 
    ANTENNAPARTIALMETALAREA 0.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
  END instr_rdata_i[19]
  PIN instr_rdata_i[18] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M3 ;
  END instr_rdata_i[18]
  PIN instr_rdata_i[17] 
    ANTENNAPARTIALMETALAREA 2.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.8559 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 173.329 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_rdata_i[17]
  PIN instr_rdata_i[16] 
    ANTENNAPARTIALMETALAREA 2.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.916 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.3423 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 124.995 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_rdata_i[16]
  PIN instr_rdata_i[15] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
  END instr_rdata_i[15]
  PIN instr_rdata_i[14] 
    ANTENNAPARTIALMETALAREA 1.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.548 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.1351 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 98.3288 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_rdata_i[14]
  PIN instr_rdata_i[13] 
    ANTENNAPARTIALMETALAREA 2.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.4189 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 99.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_rdata_i[13]
  PIN instr_rdata_i[12] 
    ANTENNAPARTIALMETALAREA 1.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.548 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.036 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 101.662 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_rdata_i[12]
  PIN instr_rdata_i[11] 
    ANTENNAPARTIALMETALAREA 2.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.991 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 119.995 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_rdata_i[11]
  PIN instr_rdata_i[10] 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.844 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.036 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 101.662 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_rdata_i[10]
  PIN instr_rdata_i[9] 
    ANTENNAPARTIALMETALAREA 1.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
  END instr_rdata_i[9]
  PIN instr_rdata_i[8] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M3 ;
  END instr_rdata_i[8]
  PIN instr_rdata_i[7] 
    ANTENNAPARTIALMETALAREA 0.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
  END instr_rdata_i[7]
  PIN instr_rdata_i[6] 
    ANTENNAPARTIALMETALAREA 1.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.66 LAYER M3 ;
  END instr_rdata_i[6]
  PIN instr_rdata_i[5] 
    ANTENNAPARTIALMETALAREA 0.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
  END instr_rdata_i[5]
  PIN instr_rdata_i[4] 
    ANTENNAPARTIALMETALAREA 1.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.66 LAYER M3 ;
  END instr_rdata_i[4]
  PIN instr_rdata_i[3] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
  END instr_rdata_i[3]
  PIN instr_rdata_i[2] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M3 ;
  END instr_rdata_i[2]
  PIN instr_rdata_i[1] 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.9685 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 96.3559 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_rdata_i[1]
  PIN instr_rdata_i[0] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.252 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.2342 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 94.9955 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_rdata_i[0]
  PIN instr_rdata_intg_i[6] 
  END instr_rdata_intg_i[6]
  PIN instr_rdata_intg_i[5] 
  END instr_rdata_intg_i[5]
  PIN instr_rdata_intg_i[4] 
  END instr_rdata_intg_i[4]
  PIN instr_rdata_intg_i[3] 
  END instr_rdata_intg_i[3]
  PIN instr_rdata_intg_i[2] 
  END instr_rdata_intg_i[2]
  PIN instr_rdata_intg_i[1] 
  END instr_rdata_intg_i[1]
  PIN instr_rdata_intg_i[0] 
  END instr_rdata_intg_i[0]
  PIN instr_err_i 
    ANTENNAPARTIALMETALAREA 2.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.14 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.8694 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 101.356 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END instr_err_i
  PIN data_req_o 
    ANTENNAPARTIALMETALAREA 1.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 41.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 153.624 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.8235 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 84.5205 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_req_o
  PIN data_gnt_i 
    ANTENNAPARTIALMETALAREA 0.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
  END data_gnt_i
  PIN data_rvalid_i 
    ANTENNAPARTIALMETALAREA 2.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M2 ;
  END data_rvalid_i
  PIN data_we_o 
    ANTENNAPARTIALMETALAREA 13.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 49.284 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 55.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 205.128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0444 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.3861 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 77.8465 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END data_we_o
  PIN data_be_o[3] 
    ANTENNAPARTIALMETALAREA 2.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 30.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 112.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.848 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.8991 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 40.3087 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0280899 LAYER VL ;
  END data_be_o[3]
  PIN data_be_o[2] 
    ANTENNAPARTIALMETALAREA 6.19 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.718 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 118.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.762 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.7412 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 32.4299 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0212653 LAYER VL ;
  END data_be_o[2]
  PIN data_be_o[1] 
    ANTENNAPARTIALMETALAREA 1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 30.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 112.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.848 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.7013 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 46.9699 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0280899 LAYER VL ;
  END data_be_o[1]
  PIN data_be_o[0] 
    ANTENNAPARTIALMETALAREA 1.15 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.07 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 31.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 115.736 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.1823 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 67.1984 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER VL ;
  END data_be_o[0]
  PIN data_addr_o[31] 
    ANTENNAPARTIALMETALAREA 0.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.1339 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 63.2705 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER VL ;
  END data_addr_o[31]
  PIN data_addr_o[30] 
    ANTENNAPARTIALMETALAREA 0.43 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.406 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.416 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4192 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.5984 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 62.1011 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END data_addr_o[30]
  PIN data_addr_o[29] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.24 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6328 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.06529 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 22.2821 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END data_addr_o[29]
  PIN data_addr_o[28] 
    ANTENNAPARTIALMETALAREA 0.27 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.016 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.9608 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.74717 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 36.0877 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END data_addr_o[28]
  PIN data_addr_o[27] 
    ANTENNAPARTIALMETALAREA 25.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 95.608 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.816 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8488 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.14396 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 21.9972 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.775194 LAYER VL ;
  END data_addr_o[27]
  PIN data_addr_o[26] 
    ANTENNAPARTIALMETALAREA 0.51 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6328 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.39498 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 31.6475 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.365621 LAYER VL ;
  END data_addr_o[26]
  PIN data_addr_o[25] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.456 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8488 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.89543 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 24.7949 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.775194 LAYER VL ;
  END data_addr_o[25]
  PIN data_addr_o[24] 
    ANTENNAPARTIALMETALAREA 23.39 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 86.358 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.616 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0736 LAYER M3 ; 
    ANTENNAMAXAREACAR 131.109 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 487.022 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER VL ;
  END data_addr_o[24]
  PIN data_addr_o[23] 
    ANTENNAPARTIALMETALAREA 24.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 88.8 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.68 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2464 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.4684 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 46.4123 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END data_addr_o[23]
  PIN data_addr_o[22] 
    ANTENNAPARTIALMETALAREA 0.43 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.406 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.784 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9184 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.75313 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 20.7322 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END data_addr_o[22]
  PIN data_addr_o[21] 
    ANTENNAPARTIALMETALAREA 21.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 80.66 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.904 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0736 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.0662 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 35.1302 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END data_addr_o[21]
  PIN data_addr_o[20] 
    ANTENNAPARTIALMETALAREA 0.59 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.152 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.0912 LAYER M3 ; 
    ANTENNAMAXAREACAR 309.449 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1144.16 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.41844 LAYER VL ;
  END data_addr_o[20]
  PIN data_addr_o[19] 
    ANTENNAPARTIALMETALAREA 0.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.152 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.53638 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 27.0545 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END data_addr_o[19]
  PIN data_addr_o[18] 
    ANTENNAPARTIALMETALAREA 16.11 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.422 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.736 LAYER M3 ; 
    ANTENNAMAXAREACAR 198.539 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 733.803 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.41844 LAYER VL ;
  END data_addr_o[18]
  PIN data_addr_o[17] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.896 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8488 LAYER M3 ; 
    ANTENNAMAXAREACAR 283.792 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1051.92 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.06383 LAYER VL ;
  END data_addr_o[17]
  PIN data_addr_o[16] 
    ANTENNAPARTIALMETALAREA 0.51 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.704 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9784 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.03185 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 32.6549 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END data_addr_o[16]
  PIN data_addr_o[15] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 119.799 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 444.315 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.634722 LAYER VL ;
  END data_addr_o[15]
  PIN data_addr_o[14] 
    ANTENNAPARTIALMETALAREA 0.43 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.406 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.408 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.12732 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 27.0824 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END data_addr_o[14]
  PIN data_addr_o[13] 
    ANTENNAPARTIALMETALAREA 13.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 51.356 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 97.976 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6328 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.70684 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 34.1152 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END data_addr_o[13]
  PIN data_addr_o[12] 
    ANTENNAPARTIALMETALAREA 15.39 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 56.758 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 29.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 111.296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.90832 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 37.4155 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END data_addr_o[12]
  PIN data_addr_o[11] 
    ANTENNAPARTIALMETALAREA 27.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 100.788 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 106.974 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 397.695 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END data_addr_o[11]
  PIN data_addr_o[10] 
    ANTENNAPARTIALMETALAREA 0.59 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 74.888 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4696 LAYER M3 ; 
    ANTENNAMAXAREACAR 168.708 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 624.899 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.775194 LAYER VL ;
  END data_addr_o[10]
  PIN data_addr_o[9] 
    ANTENNAPARTIALMETALAREA 0.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8056 LAYER M3 ; 
    ANTENNAMAXAREACAR 85.5943 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 317.372 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END data_addr_o[9]
  PIN data_addr_o[8] 
    ANTENNAPARTIALMETALAREA 14.75 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 54.39 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.864 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.7454 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 25.6693 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END data_addr_o[8]
  PIN data_addr_o[7] 
    ANTENNAPARTIALMETALAREA 13.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 49.432 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 89.392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8656 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.7318 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 81.5995 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END data_addr_o[7]
  PIN data_addr_o[6] 
    ANTENNAPARTIALMETALAREA 24.75 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 91.39 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 70.744 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2612 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.2912 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 79.2403 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.775194 LAYER VL ;
  END data_addr_o[6]
  PIN data_addr_o[5] 
    ANTENNAPARTIALMETALAREA 15.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.46 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.232 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.0245 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 116.532 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.775194 LAYER VL ;
  END data_addr_o[5]
  PIN data_addr_o[4] 
    ANTENNAPARTIALMETALAREA 0.27 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.632 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1128 LAYER M3 ; 
    ANTENNAMAXAREACAR 172.362 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 642.181 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END data_addr_o[4]
  PIN data_addr_o[3] 
    ANTENNAPARTIALMETALAREA 0.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 89.688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 9.396 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.75085 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 10.0169 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.00851426 LAYER VL ;
  END data_addr_o[3]
  PIN data_addr_o[2] 
    ANTENNAPARTIALMETALAREA 0.35 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6328 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.8969 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 43.8591 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VL ;
  END data_addr_o[2]
  PIN data_wdata_o[31] 
    ANTENNAPARTIALMETALAREA 1.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.144 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.968 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.12652 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 30.1417 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[31]
  PIN data_wdata_o[30] 
    ANTENNAPARTIALMETALAREA 2.03 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.864 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.46742 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 12.903 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[30]
  PIN data_wdata_o[29] 
    ANTENNAPARTIALMETALAREA 3.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.284 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.648 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.6303 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.80682 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[29]
  PIN data_wdata_o[28] 
    ANTENNAPARTIALMETALAREA 7.71 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.342 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.832 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.80909 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 10.4254 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[28]
  PIN data_wdata_o[27] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.536 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.78561 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 10.3803 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[27]
  PIN data_wdata_o[26] 
    ANTENNAPARTIALMETALAREA 1.23 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.366 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.11894 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.98485 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[26]
  PIN data_wdata_o[25] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.168 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.46364 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.25909 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[25]
  PIN data_wdata_o[24] 
    ANTENNAPARTIALMETALAREA 4.83 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.686 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.464 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.47879 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.24621 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[24]
  PIN data_wdata_o[23] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.208 LAYER M3 ;
  END data_wdata_o[23]
  PIN data_wdata_o[22] 
    ANTENNAPARTIALMETALAREA 1.95 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.22879 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.62121 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[22]
  PIN data_wdata_o[21] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.09621 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.20076 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[21]
  PIN data_wdata_o[20] 
    ANTENNAPARTIALMETALAREA 0.51 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.58485 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 17.0318 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[20]
  PIN data_wdata_o[19] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.929545 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.51288 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[19]
  PIN data_wdata_o[18] 
    ANTENNAPARTIALMETALAREA 0.59 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.96 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.0697 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 11.4258 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[18]
  PIN data_wdata_o[17] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.08864 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 11.5015 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[17]
  PIN data_wdata_o[16] 
    ANTENNAPARTIALMETALAREA 3.87 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.134 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.588636 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2.25152 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[16]
  PIN data_wdata_o[15] 
    ANTENNAPARTIALMETALAREA 9.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.892 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
  END data_wdata_o[15]
  PIN data_wdata_o[14] 
    ANTENNAPARTIALMETALAREA 0.59 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.15682 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.35379 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[14]
  PIN data_wdata_o[13] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.376515 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.53788 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[13]
  PIN data_wdata_o[12] 
    ANTENNAPARTIALMETALAREA 0.51 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER M3 ;
  END data_wdata_o[12]
  PIN data_wdata_o[11] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.853788 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.23258 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[11]
  PIN data_wdata_o[10] 
    ANTENNAPARTIALMETALAREA 0.59 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.328 LAYER M3 ;
  END data_wdata_o[10]
  PIN data_wdata_o[9] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.82348 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 10.5205 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[9]
  PIN data_wdata_o[8] 
    ANTENNAPARTIALMETALAREA 4.19 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.318 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.15682 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.35379 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[8]
  PIN data_wdata_o[7] 
    ANTENNAPARTIALMETALAREA 9.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.892 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.128 LAYER M3 ;
  END data_wdata_o[7]
  PIN data_wdata_o[6] 
    ANTENNAPARTIALMETALAREA 2.03 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.29318 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.55833 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[6]
  PIN data_wdata_o[5] 
    ANTENNAPARTIALMETALAREA 3.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.284 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.36 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.5697 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.88258 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[5]
  PIN data_wdata_o[4] 
    ANTENNAPARTIALMETALAREA 8.59 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.598 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.80455 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 14.1515 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[4]
  PIN data_wdata_o[3] 
    ANTENNAPARTIALMETALAREA 2.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.8197 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 10.5076 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[3]
  PIN data_wdata_o[2] 
    ANTENNAPARTIALMETALAREA 5.71 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.942 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.016 LAYER M3 ;
  END data_wdata_o[2]
  PIN data_wdata_o[1] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.536 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.60379 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 17.1076 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[1]
  PIN data_wdata_o[0] 
    ANTENNAPARTIALMETALAREA 4.27 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.614 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.384 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.23636 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 12.0492 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0378788 LAYER VL ;
  END data_wdata_o[0]
  PIN data_rdata_i[31] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
  END data_rdata_i[31]
  PIN data_rdata_i[30] 
    ANTENNAPARTIALMETALAREA 0.43 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.406 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
  END data_rdata_i[30]
  PIN data_rdata_i[29] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
  END data_rdata_i[29]
  PIN data_rdata_i[28] 
    ANTENNAPARTIALMETALAREA 2.11 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.622 LAYER M2 ;
  END data_rdata_i[28]
  PIN data_rdata_i[27] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
  END data_rdata_i[27]
  PIN data_rdata_i[26] 
    ANTENNAPARTIALMETALAREA 0.43 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.406 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.92 LAYER M3 ;
  END data_rdata_i[26]
  PIN data_rdata_i[25] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.956 LAYER M2 ;
  END data_rdata_i[25]
  PIN data_rdata_i[24] 
    ANTENNAPARTIALMETALAREA 1.95 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M2 ;
  END data_rdata_i[24]
  PIN data_rdata_i[23] 
    ANTENNAPARTIALMETALAREA 0.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
  END data_rdata_i[23]
  PIN data_rdata_i[22] 
    ANTENNAPARTIALMETALAREA 0.43 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.406 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.4414 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 119.995 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END data_rdata_i[22]
  PIN data_rdata_i[21] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.956 LAYER M2 ;
  END data_rdata_i[21]
  PIN data_rdata_i[20] 
    ANTENNAPARTIALMETALAREA 0.35 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
  END data_rdata_i[20]
  PIN data_rdata_i[19] 
    ANTENNAPARTIALMETALAREA 0.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M2 ;
  END data_rdata_i[19]
  PIN data_rdata_i[18] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.148 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.6982 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 23.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END data_rdata_i[18]
  PIN data_rdata_i[17] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
  END data_rdata_i[17]
  PIN data_rdata_i[16] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.148 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
  END data_rdata_i[16]
  PIN data_rdata_i[15] 
    ANTENNAPARTIALMETALAREA 2.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.916 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
  END data_rdata_i[15]
  PIN data_rdata_i[14] 
    ANTENNAPARTIALMETALAREA 0.59 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
  END data_rdata_i[14]
  PIN data_rdata_i[13] 
    ANTENNAPARTIALMETALAREA 0.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
  END data_rdata_i[13]
  PIN data_rdata_i[12] 
    ANTENNAPARTIALMETALAREA 0.43 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.406 LAYER M2 ;
  END data_rdata_i[12]
  PIN data_rdata_i[11] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.736 LAYER M3 ;
  END data_rdata_i[11]
  PIN data_rdata_i[10] 
    ANTENNAPARTIALMETALAREA 0.51 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M2 ;
  END data_rdata_i[10]
  PIN data_rdata_i[9] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.956 LAYER M2 ;
  END data_rdata_i[9]
  PIN data_rdata_i[8] 
    ANTENNAPARTIALMETALAREA 0.67 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.294 LAYER M2 ;
  END data_rdata_i[8]
  PIN data_rdata_i[7] 
    ANTENNAPARTIALMETALAREA 0.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M2 ;
  END data_rdata_i[7]
  PIN data_rdata_i[6] 
    ANTENNAPARTIALMETALAREA 1.95 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M2 ;
  END data_rdata_i[6]
  PIN data_rdata_i[5] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.956 LAYER M2 ;
  END data_rdata_i[5]
  PIN data_rdata_i[4] 
    ANTENNAPARTIALMETALAREA 0.27 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
  END data_rdata_i[4]
  PIN data_rdata_i[3] 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.252 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
  END data_rdata_i[3]
  PIN data_rdata_i[2] 
    ANTENNAPARTIALMETALAREA 0.35 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M2 ;
  END data_rdata_i[2]
  PIN data_rdata_i[1] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M2 ;
  END data_rdata_i[1]
  PIN data_rdata_i[0] 
    ANTENNAPARTIALMETALAREA 0.51 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M2 ;
  END data_rdata_i[0]
  PIN data_rdata_intg_i[6] 
  END data_rdata_intg_i[6]
  PIN data_rdata_intg_i[5] 
  END data_rdata_intg_i[5]
  PIN data_rdata_intg_i[4] 
  END data_rdata_intg_i[4]
  PIN data_rdata_intg_i[3] 
  END data_rdata_intg_i[3]
  PIN data_rdata_intg_i[2] 
  END data_rdata_intg_i[2]
  PIN data_rdata_intg_i[1] 
  END data_rdata_intg_i[1]
  PIN data_rdata_intg_i[0] 
  END data_rdata_intg_i[0]
  PIN data_err_i 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER M3 ;
  END data_err_i
  PIN irq_software_i 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M3 ;
  END irq_software_i
  PIN irq_timer_i 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M3 ;
  END irq_timer_i
  PIN irq_external_i 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M3 ;
  END irq_external_i
  PIN irq_fast_i[14] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M3 ;
  END irq_fast_i[14]
  PIN irq_fast_i[13] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M3 ;
  END irq_fast_i[13]
  PIN irq_fast_i[12] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1608 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.8259 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 60.2164 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.497512 LAYER VL ;
  END irq_fast_i[12]
  PIN irq_fast_i[11] 
    ANTENNAPARTIALMETALAREA 1.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.884 LAYER M3 ;
  END irq_fast_i[11]
  PIN irq_fast_i[10] 
    ANTENNAPARTIALMETALAREA 0.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1608 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.8458 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 59.6493 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.497512 LAYER VL ;
  END irq_fast_i[10]
  PIN irq_fast_i[9] 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M3 ;
  END irq_fast_i[9]
  PIN irq_fast_i[8] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1608 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.602 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 55.0473 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.497512 LAYER VL ;
  END irq_fast_i[8]
  PIN irq_fast_i[7] 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1608 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.7264 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 55.5075 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.497512 LAYER VL ;
  END irq_fast_i[7]
  PIN irq_fast_i[6] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1608 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.8507 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 55.9677 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.497512 LAYER VL ;
  END irq_fast_i[6]
  PIN irq_fast_i[5] 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M3 ;
  END irq_fast_i[5]
  PIN irq_fast_i[4] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.886 LAYER M3 ;
  END irq_fast_i[4]
  PIN irq_fast_i[3] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1608 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.1244 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 61.4851 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.497512 LAYER VL ;
  END irq_fast_i[3]
  PIN irq_fast_i[2] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M3 ;
  END irq_fast_i[2]
  PIN irq_fast_i[1] 
    ANTENNAPARTIALMETALAREA 0.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3 ;
  END irq_fast_i[1]
  PIN irq_fast_i[0] 
    ANTENNAPARTIALMETALAREA 0.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.294 LAYER M3 ;
  END irq_fast_i[0]
  PIN irq_nm_i 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1608 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.2239 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 57.3483 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.497512 LAYER VL ;
  END irq_nm_i
  PIN scramble_key_valid_i 
  END scramble_key_valid_i
  PIN scramble_key_i[127] 
  END scramble_key_i[127]
  PIN scramble_key_i[126] 
  END scramble_key_i[126]
  PIN scramble_key_i[125] 
  END scramble_key_i[125]
  PIN scramble_key_i[124] 
  END scramble_key_i[124]
  PIN scramble_key_i[123] 
  END scramble_key_i[123]
  PIN scramble_key_i[122] 
  END scramble_key_i[122]
  PIN scramble_key_i[121] 
  END scramble_key_i[121]
  PIN scramble_key_i[120] 
  END scramble_key_i[120]
  PIN scramble_key_i[119] 
  END scramble_key_i[119]
  PIN scramble_key_i[118] 
  END scramble_key_i[118]
  PIN scramble_key_i[117] 
  END scramble_key_i[117]
  PIN scramble_key_i[116] 
  END scramble_key_i[116]
  PIN scramble_key_i[115] 
  END scramble_key_i[115]
  PIN scramble_key_i[114] 
  END scramble_key_i[114]
  PIN scramble_key_i[113] 
  END scramble_key_i[113]
  PIN scramble_key_i[112] 
  END scramble_key_i[112]
  PIN scramble_key_i[111] 
  END scramble_key_i[111]
  PIN scramble_key_i[110] 
  END scramble_key_i[110]
  PIN scramble_key_i[109] 
  END scramble_key_i[109]
  PIN scramble_key_i[108] 
  END scramble_key_i[108]
  PIN scramble_key_i[107] 
  END scramble_key_i[107]
  PIN scramble_key_i[106] 
  END scramble_key_i[106]
  PIN scramble_key_i[105] 
  END scramble_key_i[105]
  PIN scramble_key_i[104] 
  END scramble_key_i[104]
  PIN scramble_key_i[103] 
  END scramble_key_i[103]
  PIN scramble_key_i[102] 
  END scramble_key_i[102]
  PIN scramble_key_i[101] 
  END scramble_key_i[101]
  PIN scramble_key_i[100] 
  END scramble_key_i[100]
  PIN scramble_key_i[99] 
  END scramble_key_i[99]
  PIN scramble_key_i[98] 
  END scramble_key_i[98]
  PIN scramble_key_i[97] 
  END scramble_key_i[97]
  PIN scramble_key_i[96] 
  END scramble_key_i[96]
  PIN scramble_key_i[95] 
  END scramble_key_i[95]
  PIN scramble_key_i[94] 
  END scramble_key_i[94]
  PIN scramble_key_i[93] 
  END scramble_key_i[93]
  PIN scramble_key_i[92] 
  END scramble_key_i[92]
  PIN scramble_key_i[91] 
  END scramble_key_i[91]
  PIN scramble_key_i[90] 
  END scramble_key_i[90]
  PIN scramble_key_i[89] 
  END scramble_key_i[89]
  PIN scramble_key_i[88] 
  END scramble_key_i[88]
  PIN scramble_key_i[87] 
  END scramble_key_i[87]
  PIN scramble_key_i[86] 
  END scramble_key_i[86]
  PIN scramble_key_i[85] 
  END scramble_key_i[85]
  PIN scramble_key_i[84] 
  END scramble_key_i[84]
  PIN scramble_key_i[83] 
  END scramble_key_i[83]
  PIN scramble_key_i[82] 
  END scramble_key_i[82]
  PIN scramble_key_i[81] 
  END scramble_key_i[81]
  PIN scramble_key_i[80] 
  END scramble_key_i[80]
  PIN scramble_key_i[79] 
  END scramble_key_i[79]
  PIN scramble_key_i[78] 
  END scramble_key_i[78]
  PIN scramble_key_i[77] 
  END scramble_key_i[77]
  PIN scramble_key_i[76] 
  END scramble_key_i[76]
  PIN scramble_key_i[75] 
  END scramble_key_i[75]
  PIN scramble_key_i[74] 
  END scramble_key_i[74]
  PIN scramble_key_i[73] 
  END scramble_key_i[73]
  PIN scramble_key_i[72] 
  END scramble_key_i[72]
  PIN scramble_key_i[71] 
  END scramble_key_i[71]
  PIN scramble_key_i[70] 
  END scramble_key_i[70]
  PIN scramble_key_i[69] 
  END scramble_key_i[69]
  PIN scramble_key_i[68] 
  END scramble_key_i[68]
  PIN scramble_key_i[67] 
  END scramble_key_i[67]
  PIN scramble_key_i[66] 
  END scramble_key_i[66]
  PIN scramble_key_i[65] 
  END scramble_key_i[65]
  PIN scramble_key_i[64] 
  END scramble_key_i[64]
  PIN scramble_key_i[63] 
  END scramble_key_i[63]
  PIN scramble_key_i[62] 
  END scramble_key_i[62]
  PIN scramble_key_i[61] 
  END scramble_key_i[61]
  PIN scramble_key_i[60] 
  END scramble_key_i[60]
  PIN scramble_key_i[59] 
  END scramble_key_i[59]
  PIN scramble_key_i[58] 
  END scramble_key_i[58]
  PIN scramble_key_i[57] 
  END scramble_key_i[57]
  PIN scramble_key_i[56] 
  END scramble_key_i[56]
  PIN scramble_key_i[55] 
  END scramble_key_i[55]
  PIN scramble_key_i[54] 
  END scramble_key_i[54]
  PIN scramble_key_i[53] 
  END scramble_key_i[53]
  PIN scramble_key_i[52] 
  END scramble_key_i[52]
  PIN scramble_key_i[51] 
  END scramble_key_i[51]
  PIN scramble_key_i[50] 
  END scramble_key_i[50]
  PIN scramble_key_i[49] 
  END scramble_key_i[49]
  PIN scramble_key_i[48] 
  END scramble_key_i[48]
  PIN scramble_key_i[47] 
  END scramble_key_i[47]
  PIN scramble_key_i[46] 
  END scramble_key_i[46]
  PIN scramble_key_i[45] 
  END scramble_key_i[45]
  PIN scramble_key_i[44] 
  END scramble_key_i[44]
  PIN scramble_key_i[43] 
  END scramble_key_i[43]
  PIN scramble_key_i[42] 
  END scramble_key_i[42]
  PIN scramble_key_i[41] 
  END scramble_key_i[41]
  PIN scramble_key_i[40] 
  END scramble_key_i[40]
  PIN scramble_key_i[39] 
  END scramble_key_i[39]
  PIN scramble_key_i[38] 
  END scramble_key_i[38]
  PIN scramble_key_i[37] 
  END scramble_key_i[37]
  PIN scramble_key_i[36] 
  END scramble_key_i[36]
  PIN scramble_key_i[35] 
  END scramble_key_i[35]
  PIN scramble_key_i[34] 
  END scramble_key_i[34]
  PIN scramble_key_i[33] 
  END scramble_key_i[33]
  PIN scramble_key_i[32] 
  END scramble_key_i[32]
  PIN scramble_key_i[31] 
  END scramble_key_i[31]
  PIN scramble_key_i[30] 
  END scramble_key_i[30]
  PIN scramble_key_i[29] 
  END scramble_key_i[29]
  PIN scramble_key_i[28] 
  END scramble_key_i[28]
  PIN scramble_key_i[27] 
  END scramble_key_i[27]
  PIN scramble_key_i[26] 
  END scramble_key_i[26]
  PIN scramble_key_i[25] 
  END scramble_key_i[25]
  PIN scramble_key_i[24] 
  END scramble_key_i[24]
  PIN scramble_key_i[23] 
  END scramble_key_i[23]
  PIN scramble_key_i[22] 
  END scramble_key_i[22]
  PIN scramble_key_i[21] 
  END scramble_key_i[21]
  PIN scramble_key_i[20] 
  END scramble_key_i[20]
  PIN scramble_key_i[19] 
  END scramble_key_i[19]
  PIN scramble_key_i[18] 
  END scramble_key_i[18]
  PIN scramble_key_i[17] 
  END scramble_key_i[17]
  PIN scramble_key_i[16] 
  END scramble_key_i[16]
  PIN scramble_key_i[15] 
  END scramble_key_i[15]
  PIN scramble_key_i[14] 
  END scramble_key_i[14]
  PIN scramble_key_i[13] 
  END scramble_key_i[13]
  PIN scramble_key_i[12] 
  END scramble_key_i[12]
  PIN scramble_key_i[11] 
  END scramble_key_i[11]
  PIN scramble_key_i[10] 
  END scramble_key_i[10]
  PIN scramble_key_i[9] 
  END scramble_key_i[9]
  PIN scramble_key_i[8] 
  END scramble_key_i[8]
  PIN scramble_key_i[7] 
  END scramble_key_i[7]
  PIN scramble_key_i[6] 
  END scramble_key_i[6]
  PIN scramble_key_i[5] 
  END scramble_key_i[5]
  PIN scramble_key_i[4] 
  END scramble_key_i[4]
  PIN scramble_key_i[3] 
  END scramble_key_i[3]
  PIN scramble_key_i[2] 
  END scramble_key_i[2]
  PIN scramble_key_i[1] 
  END scramble_key_i[1]
  PIN scramble_key_i[0] 
  END scramble_key_i[0]
  PIN scramble_nonce_i[63] 
  END scramble_nonce_i[63]
  PIN scramble_nonce_i[62] 
  END scramble_nonce_i[62]
  PIN scramble_nonce_i[61] 
  END scramble_nonce_i[61]
  PIN scramble_nonce_i[60] 
  END scramble_nonce_i[60]
  PIN scramble_nonce_i[59] 
  END scramble_nonce_i[59]
  PIN scramble_nonce_i[58] 
  END scramble_nonce_i[58]
  PIN scramble_nonce_i[57] 
  END scramble_nonce_i[57]
  PIN scramble_nonce_i[56] 
  END scramble_nonce_i[56]
  PIN scramble_nonce_i[55] 
  END scramble_nonce_i[55]
  PIN scramble_nonce_i[54] 
  END scramble_nonce_i[54]
  PIN scramble_nonce_i[53] 
  END scramble_nonce_i[53]
  PIN scramble_nonce_i[52] 
  END scramble_nonce_i[52]
  PIN scramble_nonce_i[51] 
  END scramble_nonce_i[51]
  PIN scramble_nonce_i[50] 
  END scramble_nonce_i[50]
  PIN scramble_nonce_i[49] 
  END scramble_nonce_i[49]
  PIN scramble_nonce_i[48] 
  END scramble_nonce_i[48]
  PIN scramble_nonce_i[47] 
  END scramble_nonce_i[47]
  PIN scramble_nonce_i[46] 
  END scramble_nonce_i[46]
  PIN scramble_nonce_i[45] 
  END scramble_nonce_i[45]
  PIN scramble_nonce_i[44] 
  END scramble_nonce_i[44]
  PIN scramble_nonce_i[43] 
  END scramble_nonce_i[43]
  PIN scramble_nonce_i[42] 
  END scramble_nonce_i[42]
  PIN scramble_nonce_i[41] 
  END scramble_nonce_i[41]
  PIN scramble_nonce_i[40] 
  END scramble_nonce_i[40]
  PIN scramble_nonce_i[39] 
  END scramble_nonce_i[39]
  PIN scramble_nonce_i[38] 
  END scramble_nonce_i[38]
  PIN scramble_nonce_i[37] 
  END scramble_nonce_i[37]
  PIN scramble_nonce_i[36] 
  END scramble_nonce_i[36]
  PIN scramble_nonce_i[35] 
  END scramble_nonce_i[35]
  PIN scramble_nonce_i[34] 
  END scramble_nonce_i[34]
  PIN scramble_nonce_i[33] 
  END scramble_nonce_i[33]
  PIN scramble_nonce_i[32] 
  END scramble_nonce_i[32]
  PIN scramble_nonce_i[31] 
  END scramble_nonce_i[31]
  PIN scramble_nonce_i[30] 
  END scramble_nonce_i[30]
  PIN scramble_nonce_i[29] 
  END scramble_nonce_i[29]
  PIN scramble_nonce_i[28] 
  END scramble_nonce_i[28]
  PIN scramble_nonce_i[27] 
  END scramble_nonce_i[27]
  PIN scramble_nonce_i[26] 
  END scramble_nonce_i[26]
  PIN scramble_nonce_i[25] 
  END scramble_nonce_i[25]
  PIN scramble_nonce_i[24] 
  END scramble_nonce_i[24]
  PIN scramble_nonce_i[23] 
  END scramble_nonce_i[23]
  PIN scramble_nonce_i[22] 
  END scramble_nonce_i[22]
  PIN scramble_nonce_i[21] 
  END scramble_nonce_i[21]
  PIN scramble_nonce_i[20] 
  END scramble_nonce_i[20]
  PIN scramble_nonce_i[19] 
  END scramble_nonce_i[19]
  PIN scramble_nonce_i[18] 
  END scramble_nonce_i[18]
  PIN scramble_nonce_i[17] 
  END scramble_nonce_i[17]
  PIN scramble_nonce_i[16] 
  END scramble_nonce_i[16]
  PIN scramble_nonce_i[15] 
  END scramble_nonce_i[15]
  PIN scramble_nonce_i[14] 
  END scramble_nonce_i[14]
  PIN scramble_nonce_i[13] 
  END scramble_nonce_i[13]
  PIN scramble_nonce_i[12] 
  END scramble_nonce_i[12]
  PIN scramble_nonce_i[11] 
  END scramble_nonce_i[11]
  PIN scramble_nonce_i[10] 
  END scramble_nonce_i[10]
  PIN scramble_nonce_i[9] 
  END scramble_nonce_i[9]
  PIN scramble_nonce_i[8] 
  END scramble_nonce_i[8]
  PIN scramble_nonce_i[7] 
  END scramble_nonce_i[7]
  PIN scramble_nonce_i[6] 
  END scramble_nonce_i[6]
  PIN scramble_nonce_i[5] 
  END scramble_nonce_i[5]
  PIN scramble_nonce_i[4] 
  END scramble_nonce_i[4]
  PIN scramble_nonce_i[3] 
  END scramble_nonce_i[3]
  PIN scramble_nonce_i[2] 
  END scramble_nonce_i[2]
  PIN scramble_nonce_i[1] 
  END scramble_nonce_i[1]
  PIN scramble_nonce_i[0] 
  END scramble_nonce_i[0]
  PIN debug_req_i 
    ANTENNAPARTIALMETALAREA 1.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.66 LAYER M3 ;
  END debug_req_i
  PIN crash_dump_o[159] 
    ANTENNAPARTIALMETALAREA 2.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 45.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 167.24 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5772 LAYER M3 ; 
    ANTENNAMAXAREACAR 204.82 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 759.213 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.961538 LAYER VL ;
  END crash_dump_o[159]
  PIN crash_dump_o[158] 
    ANTENNAPARTIALMETALAREA 5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.5 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 45.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 168.72 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.0552 LAYER M3 ; 
    ANTENNAMAXAREACAR 166.234 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 616.503 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[158]
  PIN crash_dump_o[157] 
    ANTENNAPARTIALMETALAREA 4.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.504 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 97.68 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8032 LAYER M3 ; 
    ANTENNAMAXAREACAR 90.1189 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 334.408 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.591693 LAYER VL ;
  END crash_dump_o[157]
  PIN crash_dump_o[156] 
    ANTENNAPARTIALMETALAREA 3.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.172 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 29.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 111 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7336 LAYER M3 ; 
    ANTENNAMAXAREACAR 397.553 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1473.06 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[156]
  PIN crash_dump_o[155] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 94.424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7144 LAYER M3 ; 
    ANTENNAMAXAREACAR 126.812 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.888 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.411523 LAYER VL ;
  END crash_dump_o[155]
  PIN crash_dump_o[154] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 70.744 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7096 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.8533 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 54.0899 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.36213 LAYER VL ;
  END crash_dump_o[154]
  PIN crash_dump_o[153] 
    ANTENNAPARTIALMETALAREA 1.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.364 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 101.528 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2756 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.9779 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 59.5146 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END crash_dump_o[153]
  PIN crash_dump_o[152] 
    ANTENNAPARTIALMETALAREA 4.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.02 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 100.936 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2756 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.8957 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 54.045 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END crash_dump_o[152]
  PIN crash_dump_o[151] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.016 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.848 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.65636 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.5037 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0280899 LAYER VL ;
  END crash_dump_o[151]
  PIN crash_dump_o[150] 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.028 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.68 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.52 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.07636 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.47205 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0227273 LAYER VL ;
  END crash_dump_o[150]
  PIN crash_dump_o[149] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 100.048 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8032 LAYER M3 ; 
    ANTENNAMAXAREACAR 102.434 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 379.974 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.591693 LAYER VL ;
  END crash_dump_o[149]
  PIN crash_dump_o[148] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 33.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 124.32 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2756 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.908 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 66.591 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END crash_dump_o[148]
  PIN crash_dump_o[147] 
    ANTENNAPARTIALMETALAREA 6.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.36 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1868 LAYER M3 ; 
    ANTENNAMAXAREACAR 63.4917 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 236.077 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[147]
  PIN crash_dump_o[146] 
    ANTENNAPARTIALMETALAREA 1.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.364 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 31.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 118.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1488 LAYER M3 ; 
    ANTENNAMAXAREACAR 113.617 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 421.165 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END crash_dump_o[146]
  PIN crash_dump_o[145] 
    ANTENNAPARTIALMETALAREA 6.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.456 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 122.248 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6088 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.8768 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 57.2038 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END crash_dump_o[145]
  PIN crash_dump_o[144] 
    ANTENNAPARTIALMETALAREA 0.92 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.404 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 80.512 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2756 LAYER M3 ; 
    ANTENNAMAXAREACAR 78.3208 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 292.043 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[144]
  PIN crash_dump_o[143] 
    ANTENNAPARTIALMETALAREA 3.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.616 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.144 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.52 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.576364 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.92205 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0227273 LAYER VL ;
  END crash_dump_o[143]
  PIN crash_dump_o[142] 
    ANTENNAPARTIALMETALAREA 2.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.324 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.52 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.667273 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2.27 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0227273 LAYER VL ;
  END crash_dump_o[142]
  PIN crash_dump_o[141] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 29.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 110.408 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2036 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.9736 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 83.4323 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END crash_dump_o[141]
  PIN crash_dump_o[140] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 36.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 136.16 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9544 LAYER M3 ; 
    ANTENNAMAXAREACAR 188.775 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 699.571 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END crash_dump_o[140]
  PIN crash_dump_o[139] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 35.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 131.424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9064 LAYER M3 ; 
    ANTENNAMAXAREACAR 175.618 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 651.233 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END crash_dump_o[139]
  PIN crash_dump_o[138] 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.028 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 39.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 148 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 70.934 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 263.041 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END crash_dump_o[138]
  PIN crash_dump_o[137] 
    ANTENNAPARTIALMETALAREA 4.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.872 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 38.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 142.08 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2756 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.5156 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 189.098 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER VL ;
  END crash_dump_o[137]
  PIN crash_dump_o[136] 
    ANTENNAPARTIALMETALAREA 1.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.292 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 35.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 132.904 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.362 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.0114 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 92.7326 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END crash_dump_o[136]
  PIN crash_dump_o[135] 
    ANTENNAPARTIALMETALAREA 2.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 36.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 134.976 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.266 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.4243 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 129.561 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END crash_dump_o[135]
  PIN crash_dump_o[134] 
    ANTENNAPARTIALMETALAREA 1.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.996 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 30.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 114.552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.362 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.3907 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 82.9737 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END crash_dump_o[134]
  PIN crash_dump_o[133] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 33.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 123.432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.266 LAYER M3 ; 
    ANTENNAMAXAREACAR 53.6801 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 198.082 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.5873 LAYER VL ;
  END crash_dump_o[133]
  PIN crash_dump_o[132] 
    ANTENNAPARTIALMETALAREA 1.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.588 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 85.248 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7792 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.1083 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 38.4557 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.724638 LAYER VL ;
  END crash_dump_o[132]
  PIN crash_dump_o[131] 
    ANTENNAPARTIALMETALAREA 0.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 77.848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.278 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.1396 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 44.3132 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.30303 LAYER VL ;
  END crash_dump_o[131]
  PIN crash_dump_o[130] 
    ANTENNAPARTIALMETALAREA 0.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 101.528 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.3984 LAYER M3 ; 
    ANTENNAMAXAREACAR 43.5958 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 161.171 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.735294 LAYER VL ;
  END crash_dump_o[130]
  PIN crash_dump_o[129] 
    ANTENNAPARTIALMETALAREA 2.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 69.56 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.7004 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.7216 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 61.7664 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.537634 LAYER VL ;
  END crash_dump_o[129]
  PIN crash_dump_o[127] 
    ANTENNAPARTIALMETALAREA 2.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.36 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 34.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 129.648 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1784 LAYER M3 ; 
    ANTENNAMAXAREACAR 74.5848 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 277.189 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[127]
  PIN crash_dump_o[126] 
    ANTENNAPARTIALMETALAREA 4.68 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.316 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.728 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1604 LAYER M3 ; 
    ANTENNAMAXAREACAR 168.481 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 626.392 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[126]
  PIN crash_dump_o[125] 
    ANTENNAPARTIALMETALAREA 4.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.688 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 81.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1872 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.0206 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 43.7584 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[125]
  PIN crash_dump_o[124] 
    ANTENNAPARTIALMETALAREA 3.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.396 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1648 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.75739 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 28.0417 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[124]
  PIN crash_dump_o[123] 
    ANTENNAPARTIALMETALAREA 3.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.208 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6812 LAYER M3 ; 
    ANTENNAMAXAREACAR 185.922 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 690.938 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[123]
  PIN crash_dump_o[122] 
    ANTENNAPARTIALMETALAREA 5.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.276 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.576 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.4105 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 45.2854 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[122]
  PIN crash_dump_o[121] 
    ANTENNAPARTIALMETALAREA 0.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.208 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6812 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.21124 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 32.6197 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[121]
  PIN crash_dump_o[120] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.744 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.79717 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 31.7619 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[120]
  PIN crash_dump_o[119] 
    ANTENNAPARTIALMETALAREA 0.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 75.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6812 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.3971 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 52.6509 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[119]
  PIN crash_dump_o[118] 
    ANTENNAPARTIALMETALAREA 2.84 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.656 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0784 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.62137 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 27.9685 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[118]
  PIN crash_dump_o[117] 
    ANTENNAPARTIALMETALAREA 8.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.044 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.544 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1872 LAYER M3 ; 
    ANTENNAMAXAREACAR 66.4001 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 245.989 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[117]
  PIN crash_dump_o[116] 
    ANTENNAPARTIALMETALAREA 2.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.212 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 67.784 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3376 LAYER M3 ; 
    ANTENNAMAXAREACAR 170.875 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 635.788 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[116]
  PIN crash_dump_o[115] 
    ANTENNAPARTIALMETALAREA 6.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.384 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6812 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.50115 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 38.8587 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[115]
  PIN crash_dump_o[114] 
    ANTENNAPARTIALMETALAREA 1.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.92 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0784 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.63288 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 27.5812 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[114]
  PIN crash_dump_o[113] 
    ANTENNAPARTIALMETALAREA 6.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.308 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 95.608 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1872 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.03054 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 36.4723 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[113]
  PIN crash_dump_o[112] 
    ANTENNAPARTIALMETALAREA 4.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.612 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.784 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3376 LAYER M3 ; 
    ANTENNAMAXAREACAR 201.2 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 748.036 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[112]
  PIN crash_dump_o[111] 
    ANTENNAPARTIALMETALAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.32 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 82.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1872 LAYER M3 ; 
    ANTENNAMAXAREACAR 77.8565 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 288.378 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[111]
  PIN crash_dump_o[110] 
    ANTENNAPARTIALMETALAREA 2.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.844 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2708 LAYER M3 ; 
    ANTENNAMAXAREACAR 170.963 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 634.818 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[110]
  PIN crash_dump_o[109] 
    ANTENNAPARTIALMETALAREA 4.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.984 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 59.496 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1872 LAYER M3 ; 
    ANTENNAMAXAREACAR 90.2743 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 334.253 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[109]
  PIN crash_dump_o[108] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.896 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2512 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.41617 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 34.2147 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[108]
  PIN crash_dump_o[107] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 98.864 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1872 LAYER M3 ; 
    ANTENNAMAXAREACAR 63.5654 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 238.139 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[107]
  PIN crash_dump_o[106] 
    ANTENNAPARTIALMETALAREA 8.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.524 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 78.736 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2512 LAYER M3 ; 
    ANTENNAMAXAREACAR 58.6581 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 217.345 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[106]
  PIN crash_dump_o[105] 
    ANTENNAPARTIALMETALAREA 0.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.928 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1872 LAYER M3 ; 
    ANTENNAMAXAREACAR 149.205 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 555.574 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[105]
  PIN crash_dump_o[104] 
    ANTENNAPARTIALMETALAREA 0.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.812 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.792 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4196 LAYER M3 ; 
    ANTENNAMAXAREACAR 165.153 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 614.621 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[104]
  PIN crash_dump_o[103] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5776 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.88222 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 14.1827 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[103]
  PIN crash_dump_o[102] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.216 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.566 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.77714 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 30.3626 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[102]
  PIN crash_dump_o[101] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.912 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5776 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.74314 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 17.4095 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[101]
  PIN crash_dump_o[100] 
    ANTENNAPARTIALMETALAREA 22.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 83.62 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2708 LAYER M2 ; 
    ANTENNAMAXAREACAR 56.8058 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 235.275 LAYER M2 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER V2 ;
  END crash_dump_o[100]
  PIN crash_dump_o[99] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.809 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 121.437 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[99]
  PIN crash_dump_o[98] 
    ANTENNAPARTIALMETALAREA 7.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.676 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8368 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.00727 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 36.2868 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END crash_dump_o[98]
  PIN crash_dump_o[97] 
    ANTENNAPARTIALMETALAREA 2.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.064 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 43.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 163.392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.3208 LAYER M3 ; 
    ANTENNAMAXAREACAR 268.938 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 998.71 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END crash_dump_o[97]
  PIN crash_dump_o[95] 
    ANTENNAPARTIALMETALAREA 15.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.608 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.344 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8176 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.69748 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 24.8571 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER VL ;
  END crash_dump_o[95]
  PIN crash_dump_o[94] 
    ANTENNAPARTIALMETALAREA 15.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 57.276 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8176 LAYER M3 ; 
    ANTENNAMAXAREACAR 95.0135 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 352.744 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[94]
  PIN crash_dump_o[93] 
    ANTENNAPARTIALMETALAREA 2.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.36 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 177.108 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 656.491 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[93]
  PIN crash_dump_o[92] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.736 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8176 LAYER M3 ; 
    ANTENNAMAXAREACAR 79.5261 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 295.518 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[92]
  PIN crash_dump_o[91] 
    ANTENNAPARTIALMETALAREA 5.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.276 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.16 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 53.1166 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 197.799 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[91]
  PIN crash_dump_o[90] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.2079 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.92 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.241772 LAYER VL ;
  END crash_dump_o[90]
  PIN crash_dump_o[89] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.976 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.93708 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 26.7275 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[89]
  PIN crash_dump_o[88] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.3545 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 91.1341 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[88]
  PIN crash_dump_o[87] 
    ANTENNAPARTIALMETALAREA 1.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.624 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.084 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.53766 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 21.7457 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[87]
  PIN crash_dump_o[86] 
    ANTENNAPARTIALMETALAREA 27.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 103.452 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.216 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.2748 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 98.3976 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER VL ;
  END crash_dump_o[86]
  PIN crash_dump_o[85] 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.328 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.136 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 191.131 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 708.337 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[85]
  PIN crash_dump_o[84] 
    ANTENNAPARTIALMETALAREA 27.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 102.268 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.488 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.26675 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.3139 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[84]
  PIN crash_dump_o[83] 
    ANTENNAPARTIALMETALAREA 28.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 105.968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.704 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.3858 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 121.019 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[83]
  PIN crash_dump_o[82] 
    ANTENNAPARTIALMETALAREA 27.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 103.156 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.968 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.31022 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 16.0208 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[82]
  PIN crash_dump_o[81] 
    ANTENNAPARTIALMETALAREA 29.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 108.632 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.112 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.2145 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 105.074 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[81]
  PIN crash_dump_o[80] 
    ANTENNAPARTIALMETALAREA 5.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.388 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.408 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.71854 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 18.6578 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[80]
  PIN crash_dump_o[79] 
    ANTENNAPARTIALMETALAREA 35.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 131.276 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.084 LAYER M2 ; 
    ANTENNAMAXAREACAR 47.2647 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 195.73 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER V2 ;
  END crash_dump_o[79]
  PIN crash_dump_o[78] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.544 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8176 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.96439 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 22.7992 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER VL ;
  END crash_dump_o[78]
  PIN crash_dump_o[77] 
    ANTENNAPARTIALMETALAREA 2.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8176 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.9435 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 100.924 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[77]
  PIN crash_dump_o[76] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8656 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.34535 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 17.2698 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[76]
  PIN crash_dump_o[75] 
    ANTENNAPARTIALMETALAREA 6.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.144 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8176 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.9393 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 40.5907 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER VL ;
  END crash_dump_o[75]
  PIN crash_dump_o[74] 
    ANTENNAPARTIALMETALAREA 6.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.644 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.084 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.4519 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 38.7773 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[74]
  PIN crash_dump_o[73] 
    ANTENNAPARTIALMETALAREA 9.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8872 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.22544 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 20.6015 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[73]
  PIN crash_dump_o[72] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.68 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.8417 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 43.9748 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[72]
  PIN crash_dump_o[71] 
    ANTENNAPARTIALMETALAREA 9.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.52 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.61759 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 22.0243 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[71]
  PIN crash_dump_o[70] 
    ANTENNAPARTIALMETALAREA 11.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 44.252 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.1417 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 37.6046 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[70]
  PIN crash_dump_o[69] 
    ANTENNAPARTIALMETALAREA 11.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 41.736 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.576 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.084 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.07635 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 23.6301 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[69]
  PIN crash_dump_o[68] 
    ANTENNAPARTIALMETALAREA 12.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 46.324 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8656 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.80273 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 26.3622 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[68]
  PIN crash_dump_o[67] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.304 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8656 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.14421 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 27.6639 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[67]
  PIN crash_dump_o[66] 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.028 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 70.448 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8416 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.29298 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 28.0075 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.537634 LAYER VL ;
  END crash_dump_o[66]
  PIN crash_dump_o[65] 
    ANTENNAPARTIALMETALAREA 8.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.784 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 56.24 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8416 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.0211 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 44.5526 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.537634 LAYER VL ;
  END crash_dump_o[65]
  PIN crash_dump_o[64] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.912 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8272 LAYER M3 ; 
    ANTENNAMAXAREACAR 138.275 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 580.359 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.365061 LAYER VL ;
  END crash_dump_o[64]
  PIN crash_dump_o[63] 
    ANTENNAPARTIALMETALAREA 7.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.416 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 28.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 104.488 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 97.6501 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 362.494 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[63]
  PIN crash_dump_o[62] 
    ANTENNAPARTIALMETALAREA 3.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.06 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 30.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 113.96 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 97.7341 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 362.871 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[62]
  PIN crash_dump_o[61] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 35.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 131.424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 122.656 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 454.979 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[61]
  PIN crash_dump_o[60] 
    ANTENNAPARTIALMETALAREA 1.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.364 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 41.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 153.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6616 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.1805 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 62.6985 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.19048 LAYER VL ;
  END crash_dump_o[60]
  PIN crash_dump_o[59] 
    ANTENNAPARTIALMETALAREA 2.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 41.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 153.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8344 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.3415 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 65.7258 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.19048 LAYER VL ;
  END crash_dump_o[59]
  PIN crash_dump_o[58] 
    ANTENNAPARTIALMETALAREA 1.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 37.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 141.192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.8496 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 46.3033 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[58]
  PIN crash_dump_o[57] 
    ANTENNAPARTIALMETALAREA 1.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 43.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 161.32 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8344 LAYER M3 ; 
    ANTENNAMAXAREACAR 155.556 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 576.75 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[57]
  PIN crash_dump_o[56] 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 40 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 148.592 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 148.361 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 550.123 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[56]
  PIN crash_dump_o[55] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 31.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 117.808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.4182 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 44.7123 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[55]
  PIN crash_dump_o[54] 
    ANTENNAPARTIALMETALAREA 1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 39.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 147.704 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.3924 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 100.042 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[54]
  PIN crash_dump_o[53] 
    ANTENNAPARTIALMETALAREA 3.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.912 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 37.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 139.12 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 124.1 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 460.358 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[53]
  PIN crash_dump_o[52] 
    ANTENNAPARTIALMETALAREA 2.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.324 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 44.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 164.28 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8344 LAYER M3 ; 
    ANTENNAMAXAREACAR 325.288 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1205.09 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.19048 LAYER VL ;
  END crash_dump_o[52]
  PIN crash_dump_o[51] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 42.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 156.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 91.0588 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 338.107 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER VL ;
  END crash_dump_o[51]
  PIN crash_dump_o[50] 
    ANTENNAPARTIALMETALAREA 1.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.996 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 36.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 136.456 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.9984 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 65.3593 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[50]
  PIN crash_dump_o[49] 
    ANTENNAPARTIALMETALAREA 5.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.424 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 30.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 112.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 203.566 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 755.586 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.15054 LAYER VL ;
  END crash_dump_o[49]
  PIN crash_dump_o[48] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 43.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 161.32 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8368 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.277 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 58.2696 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.14943 LAYER VL ;
  END crash_dump_o[48]
  PIN crash_dump_o[47] 
    ANTENNAPARTIALMETALAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.32 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 122.248 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 123.405 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 457.789 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[47]
  PIN crash_dump_o[46] 
    ANTENNAPARTIALMETALAREA 0.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 29.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 111 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8344 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.1696 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 43.7603 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.19048 LAYER VL ;
  END crash_dump_o[46]
  PIN crash_dump_o[45] 
    ANTENNAPARTIALMETALAREA 20.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 76.368 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 101.824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.342 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 40.6555 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[45]
  PIN crash_dump_o[44] 
    ANTENNAPARTIALMETALAREA 2.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.844 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 90.872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.39779 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 33.5317 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[44]
  PIN crash_dump_o[43] 
    ANTENNAPARTIALMETALAREA 4.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.504 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 31.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 117.512 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 121.807 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 450.934 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[43]
  PIN crash_dump_o[42] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 72.816 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8344 LAYER M3 ; 
    ANTENNAMAXAREACAR 55.247 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 207.276 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.19048 LAYER VL ;
  END crash_dump_o[42]
  PIN crash_dump_o[41] 
    ANTENNAPARTIALMETALAREA 2.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 80.512 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8368 LAYER M3 ; 
    ANTENNAMAXAREACAR 98.941 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 367.236 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.14943 LAYER VL ;
  END crash_dump_o[41]
  PIN crash_dump_o[40] 
    ANTENNAPARTIALMETALAREA 15.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 57.276 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.96 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.8294 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 149.721 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[40]
  PIN crash_dump_o[39] 
    ANTENNAPARTIALMETALAREA 1.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.736 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 28.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 106.264 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 94.521 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 350.954 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[39]
  PIN crash_dump_o[38] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.956 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 28.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 107.448 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7672 LAYER M3 ; 
    ANTENNAMAXAREACAR 231.494 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 858.925 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.15054 LAYER VL ;
  END crash_dump_o[38]
  PIN crash_dump_o[37] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 119.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.5298 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 45.088 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[37]
  PIN crash_dump_o[36] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 72.224 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8368 LAYER M3 ; 
    ANTENNAMAXAREACAR 200.906 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 745.786 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.72414 LAYER VL ;
  END crash_dump_o[36]
  PIN crash_dump_o[35] 
    ANTENNAPARTIALMETALAREA 1.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8928 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.6335 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 112.355 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.411523 LAYER VL ;
  END crash_dump_o[35]
  PIN crash_dump_o[34] 
    ANTENNAPARTIALMETALAREA 7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.9 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 98.864 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.94 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.8059 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 40.229 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[34]
  PIN crash_dump_o[33] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 41 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 152.44 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7672 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.5593 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 50.9328 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER VL ;
  END crash_dump_o[33]
  PIN crash_dump_o[31] 
    ANTENNAPARTIALMETALAREA 1.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.136 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.86392 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 25.4756 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[31]
  PIN crash_dump_o[30] 
    ANTENNAPARTIALMETALAREA 12.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 45.732 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 80.216 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.2057 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 157.28 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[30]
  PIN crash_dump_o[29] 
    ANTENNAPARTIALMETALAREA 11.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 41.44 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 69.56 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.70358 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 25.9223 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[29]
  PIN crash_dump_o[28] 
    ANTENNAPARTIALMETALAREA 13.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 51.06 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 89.688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.3249 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 117.021 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[28]
  PIN crash_dump_o[27] 
    ANTENNAPARTIALMETALAREA 1.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.404 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 90.28 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.66135 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 33.2462 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[27]
  PIN crash_dump_o[26] 
    ANTENNAPARTIALMETALAREA 11.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 43.068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.656 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.364 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 143.066 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[26]
  PIN crash_dump_o[25] 
    ANTENNAPARTIALMETALAREA 0.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 89.392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 106.755 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 396.154 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[25]
  PIN crash_dump_o[24] 
    ANTENNAPARTIALMETALAREA 10.68 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 39.516 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 87.024 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.42619 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 28.6237 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[24]
  PIN crash_dump_o[23] 
    ANTENNAPARTIALMETALAREA 9.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.336 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 96.2 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.11629 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 34.8493 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[23]
  PIN crash_dump_o[22] 
    ANTENNAPARTIALMETALAREA 15.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 55.796 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 79.92 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.46182 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 28.7278 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[22]
  PIN crash_dump_o[21] 
    ANTENNAPARTIALMETALAREA 9.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.816 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 70.448 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 112.787 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 418.431 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[21]
  PIN crash_dump_o[20] 
    ANTENNAPARTIALMETALAREA 10.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 37.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 74.592 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.3867 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 128.35 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[20]
  PIN crash_dump_o[19] 
    ANTENNAPARTIALMETALAREA 9.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.632 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 93.4782 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 346.989 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[19]
  PIN crash_dump_o[18] 
    ANTENNAPARTIALMETALAREA 2.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.324 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.112 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 93.5376 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 347.208 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[18]
  PIN crash_dump_o[17] 
    ANTENNAPARTIALMETALAREA 1.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 81.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 100.593 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 373.354 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[17]
  PIN crash_dump_o[16] 
    ANTENNAPARTIALMETALAREA 3.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.172 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 70.744 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 92.4384 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 343.141 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[16]
  PIN crash_dump_o[15] 
    ANTENNAPARTIALMETALAREA 6.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 85.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 60.2099 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 223.896 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[15]
  PIN crash_dump_o[14] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 86.432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.8535 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 126.417 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[14]
  PIN crash_dump_o[13] 
    ANTENNAPARTIALMETALAREA 3.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.208 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 132.884 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 495.28 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[13]
  PIN crash_dump_o[12] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 28.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 104.192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.8025 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 54.8482 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[12]
  PIN crash_dump_o[11] 
    ANTENNAPARTIALMETALAREA 1.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 96.496 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 153.255 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 570.65 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[11]
  PIN crash_dump_o[10] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 94.72 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.52 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.42523 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 27.5583 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0227273 LAYER VL ;
  END crash_dump_o[10]
  PIN crash_dump_o[9] 
    ANTENNAPARTIALMETALAREA 1.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 99.456 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 155.94 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 580.613 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[9]
  PIN crash_dump_o[8] 
    ANTENNAPARTIALMETALAREA 2.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.732 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 91.168 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.71865 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 29.7459 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[8]
  PIN crash_dump_o[7] 
    ANTENNAPARTIALMETALAREA 1.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.512 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 97.088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 60.6859 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 224.715 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END crash_dump_o[7]
  PIN crash_dump_o[6] 
    ANTENNAPARTIALMETALAREA 6.84 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.308 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 102.416 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.065 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 41.1576 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[6]
  PIN crash_dump_o[5] 
    ANTENNAPARTIALMETALAREA 0.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 28.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 106.856 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.86683 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 33.9942 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[5]
  PIN crash_dump_o[4] 
    ANTENNAPARTIALMETALAREA 6.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.532 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 101.232 LAYER M3 ;
  END crash_dump_o[4]
  PIN crash_dump_o[3] 
    ANTENNAPARTIALMETALAREA 4.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.02 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 119.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.8709 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 40.5103 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[3]
  PIN crash_dump_o[2] 
    ANTENNAPARTIALMETALAREA 7.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.676 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 94.72 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.7857 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 44.7263 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[2]
  PIN crash_dump_o[1] 
    ANTENNAPARTIALMETALAREA 5.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.536 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 28.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 105.968 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6928 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.2942 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 39.2074 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[1]
  PIN crash_dump_o[0] 
    ANTENNAPARTIALMETALAREA 1.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.996 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 102.416 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 163.671 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 608.336 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END crash_dump_o[0]
  PIN double_fault_seen_o 
    ANTENNAPARTIALMETALAREA 27.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 102.12 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 92.944 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.004 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.93758 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 36.8471 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.512821 LAYER VL ;
  END double_fault_seen_o
  PIN fetch_enable_i[3] 
  END fetch_enable_i[3]
  PIN fetch_enable_i[2] 
  END fetch_enable_i[2]
  PIN fetch_enable_i[1] 
  END fetch_enable_i[1]
  PIN fetch_enable_i[0] 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.844 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.6982 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 23.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END fetch_enable_i[0]
  PIN core_sleep_o 
    ANTENNAPARTIALMETALAREA 0.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 84.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 312.872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.264 LAYER M3 ; 
    ANTENNAMAXAREACAR 352.805 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1306.26 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.30303 LAYER VL ;
  END core_sleep_o
  PIN scan_rst_ni 
    ANTENNAPARTIALMETALAREA 0.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
  END scan_rst_ni
  PIN test_si 
    ANTENNAPARTIALMETALAREA 0.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.4444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 128.111 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END test_si
  PIN test_so 
    ANTENNAPARTIALMETALAREA 0.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.25 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.0692 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.99975 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0246154 LAYER VL ;
  END test_so
END ibex_top

END LIBRARY
