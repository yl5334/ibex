/homes/user/stud/fall23/yl5334/ibex_/ibex/APR/innovus/ibex/ibex_top.lef